** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/DIV.sch
.subckt DIV VDD OUT IN GND
*.PININFO GND:B IN:B VDD:B OUT:B
x1 VDD A[0] A[0] net2 IN GND FF
* noconn #net2
x2 VDD A[1] A[1] net3 A[0] GND FF
* noconn #net3
x3[7] VDD OUT OUT net1 A[8] GND FF
x3[6] VDD A[8] A[8] net1 A[7] GND FF
x3[5] VDD A[7] A[7] net1 A[6] GND FF
x3[4] VDD A[6] A[6] net1 A[5] GND FF
x3[3] VDD A[5] A[5] net1 A[4] GND FF
x3[2] VDD A[4] A[4] net1 A[3] GND FF
x3[1] VDD A[3] A[3] net1 A[2] GND FF
x3[0] VDD A[2] A[2] net1 A[1] GND FF
* noconn #net1
.ends

* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/DIV/FF/FF.sym # of pins=6
** sym_path: /foss/designs/RO_Aging_UNICASS/DIV/FF/FF.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/FF/FF.sch
.subckt FF VDD D Q_N Q CLK GND
*.PININFO GND:B CLK:B VDD:B Q:B Q_N:B D:B
x1 CLKN VDD net1 D GND CLK passgate_DIV
x2 VDD net2 net1 GND inv_DIV
x3 CLK VDD net1 net4 GND CLKN passgate_DIV
x4 VDD net4 net2 GND inv_DIV
x5 CLK VDD net3 net2 GND CLKN passgate_DIV
x6 VDD net5 net3 GND inv_DIV
x7 CLKN VDD net3 Q_N GND CLK passgate_DIV
x8 VDD Q Q_N GND inv_DIV
x10 VDD CLKN CLK GND inv_DIV
x9 VDD Q_N net5 GND inv_DIV
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/DIV/passgate_DIV/passgate_DIV.sym # of pins=6
** sym_path: /foss/designs/RO_Aging_UNICASS/DIV/passgate_DIV/passgate_DIV.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/passgate_DIV/passgate_DIV.sch
.subckt passgate_DIV CLKN VDD OUT IN GND CLK
*.PININFO VDD:B OUT:B GND:B IN:B CLKN:B CLK:B
M3 IN CLK OUT GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
M1 IN CLKN OUT VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  inv_DIV.sym # of pins=4
** sym_path: /foss/designs/RO_Aging_UNICASS/DIV/inv_DIV/inv_DIV.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/inv_DIV/inv_DIV.sch
.subckt inv_DIV VDD OUT IN GND
*.PININFO VDD:B OUT:B GND:B IN:B
M3 OUT IN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
M1 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends

.end
