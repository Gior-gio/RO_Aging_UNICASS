* Extracted by KLayout with SKY130 LVS runset on : 09/11/2024 16:52

.SUBCKT FF CLK GND Q D Q_N VDD
M$1 VDD Q_N Q VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000 AS=600000000000
+ AD=600000000000 PS=5200000 PD=5200000
M$2 VDD CLK \$2 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000 AS=600000000000
+ AD=600000000000 PS=5200000 PD=5200000
M$3 VDD \$14 \$8 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000 AS=600000000000
+ AD=600000000000 PS=5200000 PD=5200000
M$4 \$20 \$2 \$21 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$6 \$14 \$13 VDD VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$9 \$15 CLK \$16 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$10 \$23 \$19 VDD VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$11 D \$2 \$12 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$13 \$17 CLK \$18 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$15 \$9 \$23 VDD VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$17 GND \$14 \$8 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$18 GND \$13 \$14 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$19 GND CLK \$2 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$20 \$20 CLK \$21 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$21 GND Q_N Q GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$22 GND \$23 \$9 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$23 GND \$19 \$23 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$24 D CLK \$12 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000 AS=195000000000
+ AD=195000000000 PS=1900000 PD=1900000
M$25 \$15 \$2 \$16 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$26 \$17 \$2 \$18 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
.ENDS FF
