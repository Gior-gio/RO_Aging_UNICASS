* Extracted by KLayout with SKY130 LVS runset on : 05/11/2024 15:06

.SUBCKT rovcel2 VSS Out IN VDD P
M$1 VDD P \$22 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=190000000
+ AS=6.25575e+13 AD=6.25575e+13 PS=221090000 PD=221090000
M$41 \$22 IN Out VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$45 Out IN VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
.ENDS rovcel2
