* Extracted by KLayout with SKY130 LVS runset on : 04/11/2024 04:09

.SUBCKT rovcel2_LVT GND OUT IN VDD
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000 AS=4.275e+12
+ AD=4.275e+12 PS=30300000 PD=30300000
M$5 OUT IN GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000 AS=1.26e+12
+ AD=1.26e+12 PS=9600000 PD=9600000
M$7 OUT GND \$28 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$8 OUT GND \$25 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$9 OUT VDD \$25 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$10 OUT VDD \$28 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
.ENDS rovcel2_LVT
