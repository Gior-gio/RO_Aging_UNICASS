magic
tech sky130
timestamp 1729529908
<< checkpaint >>
rect 0 -1 1 1
<< l67d20 >>
<< l68d20 >>
rect 0 0 1 1
<< l67d44 >>
<< l65d20 >>
rect 0 0 1 1
<< l66d44 >>
<< l66d20 >>
rect 0 -1 1 0
<< l95d20 >>
rect 0 -1 1 0
<< l65d44 >>
<< l94d20 >>
rect 0 0 1 1
<< l93d44 >>
<< l64d20 >>
rect 0 -1 1 1
<< end >>
