** sch_path: /foss/designs/RO_Aging_UNICASS/HVT/RingStage/RingStage2.sch
**.subckt RingStage2 In Out VDD VSS
*.iopin In
*.iopin Out
*.iopin VDD
*.iopin VSS
x1 VDD Out In VSS inverter
x2 Out VDD VSS VDD VSS net2 passGate_hvt
x3 Out VDD VSS VDD VSS net1 passGate_hvt
**.ends

* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/HVT/inverter/inverter.sym # of pins=4
** sym_path: /foss/designs/RO_Aging_UNICASS/HVT/inverter/inverter.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/HVT/inverter/inverter.sch
.subckt inverter VDD Out In VSS
*.iopin VDD
*.iopin Out
*.iopin VSS
*.iopin In
XM2 Out In VDD VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Out In VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/HVT/passGate_hvt/passGate_hvt.sym # of pins=6
** sym_path: /foss/designs/RO_Aging_UNICASS/HVT/passGate_hvt/passGate_hvt.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/HVT/passGate_hvt/passGate_hvt.sch
.subckt passGate_hvt In CLKN VSS VDD CLK Out
*.iopin In
*.iopin CLKN
*.iopin Out
*.iopin VSS
*.iopin VDD
*.iopin CLK
XM2 Out CLKN In VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Out CLK In VSS sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
