* Extracted by KLayout with SKY130 LVS runset on : 09/11/2024 11:56

.SUBCKT passgate_DIV GND CLK IN OUT VDD CLKN
M$1 IN CLKN OUT VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$2 IN CLK OUT GND sky130_fd_pr__nfet_01v8 L=150000 W=650000 AS=195000000000
+ AD=195000000000 PS=1900000 PD=1900000
.ENDS passgate_DIV
