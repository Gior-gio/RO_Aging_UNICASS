* Extracted by KLayout with SKY130 LVS runset on : 09/11/2024 17:04

.SUBCKT inv_DIV GND OUT IN VDD
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000 AS=600000000000
+ AD=600000000000 PS=5200000 PD=5200000
M$3 GND IN OUT GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
.ENDS inv_DIV
