* Extracted by KLayout with SKY130 LVS runset on : 10/11/2024 15:58

.SUBCKT RO_LVT_13St_x1 DUT_Gate RON Drain_Force GND Drain_Sense RO DUT_Header
+ DUT_Footer VDD OUT
M$1 \$30 \$61 \$6 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$5 VDD RON \$30 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$45 \$32 \$6 \$18 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$49 VDD DUT_Footer \$32 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$89 \$33 \$18 \$21 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$93 VDD RON \$33 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$133 \$72 VDD \$61 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$134 \$73 VDD \$61 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$135 VDD \$76 \$61 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$139 \$74 VDD \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$140 \$75 VDD \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$141 VDD \$64 \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$145 \$77 VDD \$64 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$146 \$78 VDD \$64 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$147 VDD \$81 \$64 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$151 \$6 RO DUT_Gate VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$152 \$79 VDD \$81 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$153 \$6 RO \$17 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$154 \$80 VDD \$81 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$155 VDD \$84 \$81 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$159 \$82 VDD \$84 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$160 \$83 VDD \$84 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$161 VDD \$87 \$84 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$165 \$85 VDD \$87 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$166 \$86 VDD \$87 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$167 VDD \$90 \$87 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$171 \$88 VDD \$90 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$172 \$89 VDD \$90 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$173 Drain_Force RO \$18 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=1900000
+ AS=570000000000 AD=570000000000 PS=4400000 PD=4400000
M$174 VDD \$93 \$90 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$176 Drain_Sense RO \$18 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=1900000
+ AS=570000000000 AD=570000000000 PS=4400000 PD=4400000
M$179 \$91 VDD \$93 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$180 \$92 VDD \$93 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$181 VDD \$96 \$93 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$185 \$94 VDD \$96 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$186 \$95 VDD \$96 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$187 VDD OUT \$96 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$191 \$97 VDD OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$192 \$98 VDD OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$193 VDD \$21 OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$197 \$21 VDD GND VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$198 \$21 VDD \$22 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$199 \$6 \$61 \$7 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.533e+12 AD=1.533e+12 PS=7760000 PD=7760000
M$201 \$7 RO GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.4385e+13 AD=1.4385e+13 PS=76700000 PD=76700000
M$221 \$18 \$6 \$19 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.533e+12 AD=1.533e+12 PS=7760000 PD=7760000
M$223 \$19 DUT_Header GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.4385e+13 AD=1.4385e+13 PS=76700000 PD=76700000
M$243 \$21 \$18 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.533e+12 AD=1.533e+12 PS=7760000 PD=7760000
M$245 \$72 GND \$61 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$246 \$73 GND \$61 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$247 \$61 \$76 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$249 \$74 GND \$76 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$250 \$75 GND \$76 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$251 \$76 \$64 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$253 \$77 GND \$64 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$254 \$78 GND \$64 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$255 \$64 \$81 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$257 \$6 RON DUT_Gate GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$258 \$79 GND \$81 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$259 \$6 RON \$17 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$260 \$80 GND \$81 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$261 \$81 \$84 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$263 \$82 GND \$84 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$264 \$83 GND \$84 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$265 \$84 \$87 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$267 \$85 GND \$87 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$268 \$86 GND \$87 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$269 \$87 \$90 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$271 \$88 GND \$90 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$272 \$89 GND \$90 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$273 Drain_Force RON \$18 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=420000
+ AS=126000000000 AD=126000000000 PS=1440000 PD=1440000
M$274 \$90 \$93 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$276 Drain_Sense RON \$18 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=420000
+ AS=126000000000 AD=126000000000 PS=1440000 PD=1440000
M$277 \$91 GND \$93 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$278 \$92 GND \$93 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$279 \$93 \$96 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$281 \$94 GND \$96 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$282 \$95 GND \$96 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$283 \$96 OUT GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$285 \$97 GND OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$286 \$98 GND OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$287 OUT \$21 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$289 \$21 RON GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$290 \$21 RON \$22 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
.ENDS RO_LVT_13St_x1
