** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/inv_DIV/inv_DIV.sch
.subckt inv_DIV VDD OUT IN GND
*.PININFO VDD:B OUT:B GND:B IN:B
M3 OUT IN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
M1 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=2
.ends
.end
