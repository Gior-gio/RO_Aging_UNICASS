* Extracted by KLayout with SKY130 LVS runset on : 06/11/2024 23:04

.SUBCKT rovcel1_x1_LVT GND DUT_Footer DUT_Header RO Drain_Force RON Drain_Sense
+ OUT IN VDD
M$1 \$75 IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$5 VDD DUT_Footer \$75 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$45 Drain_Force RO OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=1900000
+ AS=570000000000 AD=570000000000 PS=4400000 PD=4400000
M$46 Drain_Sense RO OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=1900000
+ AS=570000000000 AD=570000000000 PS=4400000 PD=4400000
M$47 Drain_Force RON OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=420000
+ AS=126000000000 AD=126000000000 PS=1440000 PD=1440000
M$48 Drain_Sense RON OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=420000
+ AS=126000000000 AD=126000000000 PS=1440000 PD=1440000
M$49 GND DUT_Header \$38 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.26e+13 AD=1.26e+13 PS=96000000 PD=96000000
M$69 \$38 IN OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000 AS=1.26e+12
+ AD=1.26e+12 PS=9600000 PD=9600000
.ENDS rovcel1_x1_LVT
