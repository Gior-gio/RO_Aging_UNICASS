* Extracted by KLayout with SKY130 LVS runset on : 04/11/2024 15:09

.SUBCKT MUX S[0] VSS In[11] VDD S[3] S[1] In[10] Out In[9] In[8] S[2] In[7]
+ In[6] In[5] In[4] In[3] In[2] In[1] In[0]
X$1 VSS S[0] \$7 In[11] VDD \$6 MUX_TG
X$4 VSS \$6 \$120 In[2] VDD S[0] MUX_TG
X$5 VSS \$6 \$25 In[8] VDD S[0] MUX_TG
X$6 VSS \$6 \$83 In[4] VDD S[0] MUX_TG
X$7 VSS \$6 \$139 In[0] VDD S[0] MUX_TG
X$8 VSS \$6 \$7 In[10] VDD S[0] MUX_TG
X$9 VSS \$6 \$65 In[6] VDD S[0] MUX_TG
X$33 VSS S[0] \$65 In[7] VDD \$6 MUX_TG
X$34 VSS S[0] \$25 In[9] VDD \$6 MUX_TG
X$35 VSS S[0] \$83 In[5] VDD \$6 MUX_TG
X$36 VSS S[0] \$120 In[3] VDD \$6 MUX_TG
X$37 VSS S[0] \$139 In[1] VDD \$6 MUX_TG
X$42 VSS S[1] \$132 \$120 VDD \$24 MUX_TG
X$43 VSS S[1] \$19 \$7 VDD \$24 MUX_TG
X$44 VSS \$27 \$18 \$19 VDD S[2] MUX_TG
X$45 VSS \$24 \$132 \$139 VDD S[1] MUX_TG
X$46 VSS S[2] \$96 \$81 VDD \$27 MUX_TG
X$47 VSS \$24 \$19 \$25 VDD S[1] MUX_TG
X$48 VSS \$24 \$81 \$83 VDD S[1] MUX_TG
X$49 VSS \$27 \$96 \$132 VDD S[2] MUX_TG
X$50 VSS S[3] Out \$18 VDD \$15 MUX_TG
X$51 VSS S[1] \$81 \$65 VDD \$24 MUX_TG
X$52 VSS \$15 Out \$96 VDD S[3] MUX_TG
M$1 VDD S[0] \$6 VDD sky130_fd_pr__pfet_01v8 L=150000 W=19000000 AS=6.1275e+12
+ AD=6.1275e+12 PS=26330000 PD=26330000
M$5 \$6 S[0] VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
M$7 VDD S[3] \$15 VDD sky130_fd_pr__pfet_01v8 L=150000 W=19000000 AS=6.1275e+12
+ AD=6.1275e+12 PS=26330000 PD=26330000
M$11 \$15 S[3] VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
M$13 VDD S[2] \$27 VDD sky130_fd_pr__pfet_01v8 L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$17 \$27 S[2] VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
M$19 VDD S[1] \$24 VDD sky130_fd_pr__pfet_01v8 L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$23 \$24 S[1] VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
.ENDS MUX

.SUBCKT MUX_TG VSS A Out In VDD AB
M$1 In AB Out VDD sky130_fd_pr__pfet_01v8 L=150000 W=19000000 AS=6.1275e+12
+ AD=6.1275e+12 PS=26330000 PD=26330000
M$5 Out A In VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
.ENDS MUX_TG
