* Extracted by KLayout with SKY130 LVS runset on : 07/11/2024 15:30

.SUBCKT pmos_lvt VSS VG VS VD
M$1 VS VG VD VSS sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000 AS=4.275e+12
+ AD=4.275e+12 PS=30300000 PD=30300000
.ENDS pmos_lvt
