* Extracted by KLayout with SKY130 LVS runset on : 15/10/2024 02:16

.SUBCKT TOP
X$1 OUT CLK GND IN sky130_gnd nfet$1
X$2 VDD OUT CLKN IN pfet$1
.ENDS TOP

.SUBCKT pfet$1 \$1 \$2 \$3 \$4
M$1 \$4 \$3 \$2 \$1 sky130_fd_pr__pfet_01v8 L=0.15 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$1

.SUBCKT nfet$1 \$1 \$2 \$3 \$4 sky130_gnd
M$1 \$4 \$2 \$1 sky130_gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$1
