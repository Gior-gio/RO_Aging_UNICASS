* NGSPICE file created from inverter.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_4A3DHF a_n33_n133# a_15_n45# a_n175_n219# a_n73_n45#
X0 a_15_n45# a_n33_n133# a_n73_n45# a_n175_n219# sky130_fd_pr__nfet_01v8 ad=0.1305 pd=1.48 as=0.1305 ps=1.48 w=0.45 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_hvt_HVTLRR w_n211_n309# a_15_n90# a_n33_n187# a_n73_n90#
X0 a_15_n90# a_n33_n187# a_n73_n90# w_n211_n309# sky130_fd_pr__pfet_01v8_hvt ad=0.261 pd=2.38 as=0.261 ps=2.38 w=0.9 l=0.15
.ends

.subckt inverter VDD Out In VSS
XXM1 In Out VSS VSS sky130_fd_pr__nfet_01v8_4A3DHF
XXM2 VDD Out In VDD sky130_fd_pr__pfet_01v8_hvt_HVTLRR
.ends

