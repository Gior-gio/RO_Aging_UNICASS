* Extracted by KLayout with SKY130 LVS runset on : 07/11/2024 01:09

.SUBCKT RO_LVT_13St_x1 DUT_Gate RON Drain_Force GND Drain_Sense RO DUT_Header
+ DUT_Footer VDD OUT
M$1 \$31 \$24 \$25 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$5 VDD RON \$31 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$45 \$33 \$25 \$17 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$49 VDD DUT_Footer \$33 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$89 \$34 \$17 \$26 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$93 VDD RON \$34 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$133 \$80 VDD \$24 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$134 \$81 VDD \$24 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$135 VDD \$71 \$24 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$139 \$82 VDD \$71 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$140 \$83 VDD \$71 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$141 VDD \$72 \$71 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$145 \$84 VDD \$72 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$146 \$85 VDD \$72 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$147 VDD \$73 \$72 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$151 \$25 RO DUT_Gate VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$152 \$86 VDD \$73 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$153 \$25 RO \$16 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$154 \$87 VDD \$73 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$155 VDD \$74 \$73 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$159 \$88 VDD \$74 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$160 \$89 VDD \$74 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$161 VDD \$75 \$74 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$165 \$90 VDD \$75 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$166 \$91 VDD \$75 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$167 VDD \$76 \$75 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$171 \$92 VDD \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$172 \$93 VDD \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$173 Drain_Force RO \$17 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=1900000
+ AS=570000000000 AD=570000000000 PS=4400000 PD=4400000
M$174 VDD \$77 \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$176 Drain_Sense RO \$17 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=1900000
+ AS=570000000000 AD=570000000000 PS=4400000 PD=4400000
M$179 \$94 VDD \$77 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$180 \$95 VDD \$77 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$181 VDD \$78 \$77 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$185 \$96 VDD \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$186 \$97 VDD \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$187 VDD OUT \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$191 \$98 VDD OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$192 \$99 VDD OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$193 VDD \$26 OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$197 \$26 VDD GND VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$198 \$26 VDD \$20 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$199 \$25 \$24 \$6 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$201 \$6 RO GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.26e+13 AD=1.26e+13 PS=96000000 PD=96000000
M$221 \$17 \$25 \$18 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$223 \$18 DUT_Header GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.26e+13 AD=1.26e+13 PS=96000000 PD=96000000
M$243 \$26 \$17 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$245 \$80 GND \$24 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$246 \$81 GND \$24 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$247 \$24 \$71 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$249 \$82 GND \$71 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$250 \$83 GND \$71 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$251 \$71 \$72 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$253 \$84 GND \$72 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$254 \$85 GND \$72 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$255 \$72 \$73 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$257 \$25 RON DUT_Gate GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$258 \$86 GND \$73 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$259 \$25 RON \$16 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$260 \$87 GND \$73 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$261 \$73 \$74 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$263 \$88 GND \$74 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$264 \$89 GND \$74 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$265 \$74 \$75 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$267 \$90 GND \$75 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$268 \$91 GND \$75 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$269 \$75 \$76 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$271 \$92 GND \$76 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$272 \$93 GND \$76 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$273 Drain_Force RON \$17 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=420000
+ AS=126000000000 AD=126000000000 PS=1440000 PD=1440000
M$274 \$76 \$77 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$275 Drain_Sense RON \$17 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=420000
+ AS=126000000000 AD=126000000000 PS=1440000 PD=1440000
M$277 \$94 GND \$77 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$278 \$95 GND \$77 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$279 \$77 \$78 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$281 \$96 GND \$78 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$282 \$97 GND \$78 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$283 \$78 OUT GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$285 \$98 GND OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$286 \$99 GND OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$287 OUT \$26 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$289 \$26 RON GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$290 \$26 RON \$20 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
.ENDS RO_LVT_13St_x1
