magic
tech sky130A
magscale 1 2
timestamp 1728247509
<< checkpaint >>
rect -944 -3454 2094 -3136
rect -944 -4254 4509 -3454
rect -944 -4625 323635 -4254
rect -944 -4678 326218 -4625
rect -944 -4731 326587 -4678
rect -944 -4784 326956 -4731
rect -944 -4837 327325 -4784
rect -944 -7284 327694 -4837
rect 323276 -7655 327694 -7284
rect 323645 -7708 327694 -7655
rect 324014 -7761 327694 -7708
rect 324383 -7814 327694 -7761
rect 324752 -7867 327694 -7814
<< error_s >>
rect 1505 -3821 1759 -3787
rect 1520 -3855 1539 -3842
rect 1517 -3883 1539 -3855
rect 1409 -3973 1539 -3883
rect 1725 -3855 1744 -3842
rect 1725 -3883 1747 -3855
rect 1551 -3923 1713 -3889
rect 1569 -3973 1695 -3962
rect 1725 -3973 1855 -3883
rect 1409 -4033 1855 -3973
rect 1409 -4123 1539 -4033
rect 1551 -4117 1713 -4083
rect 1517 -4151 1539 -4123
rect 1725 -4123 1855 -4033
rect 1725 -4151 1747 -4123
rect 1505 -4219 1759 -4185
rect 4066 -4207 4124 -4201
rect 4066 -4241 4078 -4207
rect 4066 -4247 4124 -4241
rect 79 -4305 333 -4271
rect 103 -4339 113 -4335
rect 91 -4367 113 -4339
rect -17 -4466 113 -4367
rect 299 -4339 309 -4335
rect 299 -4367 321 -4339
rect 125 -4407 287 -4373
rect 299 -4396 429 -4367
rect 299 -4432 465 -4396
rect 4066 -4401 4124 -4395
rect 143 -4466 269 -4455
rect 299 -4466 702 -4432
rect 4066 -4435 4078 -4401
rect 4066 -4441 4124 -4435
rect -17 -4487 465 -4466
rect -17 -4600 482 -4487
rect 668 -4500 687 -4487
rect 668 -4528 690 -4500
rect 494 -4568 656 -4534
rect 498 -4574 518 -4572
rect -17 -4602 490 -4600
rect -17 -4618 482 -4602
rect 512 -4618 638 -4607
rect 668 -4618 798 -4528
rect -17 -4622 798 -4618
rect -17 -4721 113 -4622
rect 125 -4715 287 -4681
rect 299 -4684 798 -4622
rect 299 -4700 482 -4684
rect 91 -4749 113 -4721
rect 299 -4749 490 -4700
rect 498 -4734 518 -4728
rect 316 -4783 490 -4749
rect 494 -4768 656 -4734
rect 498 -4774 518 -4768
rect 668 -4774 798 -4684
rect 2810 -4714 2844 -4696
rect 2810 -4750 2880 -4714
rect 79 -4800 490 -4783
rect 79 -4802 482 -4800
rect 668 -4802 690 -4774
rect 2827 -4784 2898 -4750
rect 79 -4817 465 -4802
rect 316 -4836 465 -4817
rect 316 -4853 702 -4836
rect 448 -4870 702 -4853
rect 1555 -5007 1613 -5001
rect 1555 -5041 1567 -5007
rect 1555 -5047 1613 -5041
rect 2827 -5135 2897 -4784
rect 3009 -4852 3067 -4846
rect 3009 -4886 3021 -4852
rect 3009 -4892 3067 -4886
rect 3203 -4905 3213 -4851
rect 3009 -5052 3067 -5046
rect 3009 -5086 3021 -5052
rect 3009 -5092 3067 -5086
rect 176 -5195 527 -5161
rect 2827 -5171 2880 -5135
rect 3257 -5188 3267 -4905
rect 3403 -5007 3461 -5001
rect 5251 -5007 5309 -5001
rect 7099 -5007 7157 -5001
rect 8947 -5007 9005 -5001
rect 10795 -5007 10853 -5001
rect 12643 -5007 12701 -5001
rect 14491 -5007 14549 -5001
rect 16339 -5007 16397 -5001
rect 18187 -5007 18245 -5001
rect 20035 -5007 20093 -5001
rect 21883 -5007 21941 -5001
rect 23731 -5007 23789 -5001
rect 25579 -5007 25637 -5001
rect 27427 -5007 27485 -5001
rect 29275 -5007 29333 -5001
rect 31123 -5007 31181 -5001
rect 32971 -5007 33029 -5001
rect 34819 -5007 34877 -5001
rect 36667 -5007 36725 -5001
rect 38515 -5007 38573 -5001
rect 40363 -5007 40421 -5001
rect 42211 -5007 42269 -5001
rect 44059 -5007 44117 -5001
rect 45907 -5007 45965 -5001
rect 47755 -5007 47813 -5001
rect 49603 -5007 49661 -5001
rect 51451 -5007 51509 -5001
rect 53299 -5007 53357 -5001
rect 55147 -5007 55205 -5001
rect 56995 -5007 57053 -5001
rect 58843 -5007 58901 -5001
rect 60691 -5007 60749 -5001
rect 62539 -5007 62597 -5001
rect 64387 -5007 64445 -5001
rect 66235 -5007 66293 -5001
rect 68083 -5007 68141 -5001
rect 69931 -5007 69989 -5001
rect 71779 -5007 71837 -5001
rect 73627 -5007 73685 -5001
rect 75475 -5007 75533 -5001
rect 77323 -5007 77381 -5001
rect 79171 -5007 79229 -5001
rect 81019 -5007 81077 -5001
rect 82867 -5007 82925 -5001
rect 84715 -5007 84773 -5001
rect 86563 -5007 86621 -5001
rect 88411 -5007 88469 -5001
rect 90259 -5007 90317 -5001
rect 92107 -5007 92165 -5001
rect 93955 -5007 94013 -5001
rect 95803 -5007 95861 -5001
rect 97651 -5007 97709 -5001
rect 99499 -5007 99557 -5001
rect 101347 -5007 101405 -5001
rect 103195 -5007 103253 -5001
rect 105043 -5007 105101 -5001
rect 106891 -5007 106949 -5001
rect 108739 -5007 108797 -5001
rect 110587 -5007 110645 -5001
rect 112435 -5007 112493 -5001
rect 114283 -5007 114341 -5001
rect 116131 -5007 116189 -5001
rect 117979 -5007 118037 -5001
rect 119827 -5007 119885 -5001
rect 121675 -5007 121733 -5001
rect 123523 -5007 123581 -5001
rect 125371 -5007 125429 -5001
rect 127219 -5007 127277 -5001
rect 129067 -5007 129125 -5001
rect 130915 -5007 130973 -5001
rect 132763 -5007 132821 -5001
rect 134611 -5007 134669 -5001
rect 136459 -5007 136517 -5001
rect 138307 -5007 138365 -5001
rect 140155 -5007 140213 -5001
rect 142003 -5007 142061 -5001
rect 143851 -5007 143909 -5001
rect 145699 -5007 145757 -5001
rect 147547 -5007 147605 -5001
rect 149395 -5007 149453 -5001
rect 151243 -5007 151301 -5001
rect 153091 -5007 153149 -5001
rect 154939 -5007 154997 -5001
rect 156787 -5007 156845 -5001
rect 158635 -5007 158693 -5001
rect 160483 -5007 160541 -5001
rect 162331 -5007 162389 -5001
rect 164179 -5007 164237 -5001
rect 166027 -5007 166085 -5001
rect 167875 -5007 167933 -5001
rect 169723 -5007 169781 -5001
rect 171571 -5007 171629 -5001
rect 173419 -5007 173477 -5001
rect 175267 -5007 175325 -5001
rect 177115 -5007 177173 -5001
rect 178963 -5007 179021 -5001
rect 3403 -5041 3415 -5007
rect 5251 -5041 5263 -5007
rect 7099 -5041 7111 -5007
rect 8947 -5041 8959 -5007
rect 10795 -5041 10807 -5007
rect 12643 -5041 12655 -5007
rect 14491 -5041 14503 -5007
rect 16339 -5041 16351 -5007
rect 18187 -5041 18199 -5007
rect 20035 -5041 20047 -5007
rect 21883 -5041 21895 -5007
rect 23731 -5041 23743 -5007
rect 25579 -5041 25591 -5007
rect 27427 -5041 27439 -5007
rect 29275 -5041 29287 -5007
rect 31123 -5041 31135 -5007
rect 32971 -5041 32983 -5007
rect 34819 -5041 34831 -5007
rect 36667 -5041 36679 -5007
rect 38515 -5041 38527 -5007
rect 40363 -5041 40375 -5007
rect 42211 -5041 42223 -5007
rect 44059 -5041 44071 -5007
rect 45907 -5041 45919 -5007
rect 47755 -5041 47767 -5007
rect 49603 -5041 49615 -5007
rect 51451 -5041 51463 -5007
rect 53299 -5041 53311 -5007
rect 55147 -5041 55159 -5007
rect 56995 -5041 57007 -5007
rect 58843 -5041 58855 -5007
rect 60691 -5041 60703 -5007
rect 62539 -5041 62551 -5007
rect 64387 -5041 64399 -5007
rect 66235 -5041 66247 -5007
rect 68083 -5041 68095 -5007
rect 69931 -5041 69943 -5007
rect 71779 -5041 71791 -5007
rect 73627 -5041 73639 -5007
rect 75475 -5041 75487 -5007
rect 77323 -5041 77335 -5007
rect 79171 -5041 79183 -5007
rect 81019 -5041 81031 -5007
rect 82867 -5041 82879 -5007
rect 84715 -5041 84727 -5007
rect 86563 -5041 86575 -5007
rect 88411 -5041 88423 -5007
rect 90259 -5041 90271 -5007
rect 92107 -5041 92119 -5007
rect 93955 -5041 93967 -5007
rect 95803 -5041 95815 -5007
rect 97651 -5041 97663 -5007
rect 99499 -5041 99511 -5007
rect 101347 -5041 101359 -5007
rect 103195 -5041 103207 -5007
rect 105043 -5041 105055 -5007
rect 106891 -5041 106903 -5007
rect 108739 -5041 108751 -5007
rect 110587 -5041 110599 -5007
rect 112435 -5041 112447 -5007
rect 114283 -5041 114295 -5007
rect 116131 -5041 116143 -5007
rect 117979 -5041 117991 -5007
rect 119827 -5041 119839 -5007
rect 121675 -5041 121687 -5007
rect 123523 -5041 123535 -5007
rect 125371 -5041 125383 -5007
rect 127219 -5041 127231 -5007
rect 129067 -5041 129079 -5007
rect 130915 -5041 130927 -5007
rect 132763 -5041 132775 -5007
rect 134611 -5041 134623 -5007
rect 136459 -5041 136471 -5007
rect 138307 -5041 138319 -5007
rect 140155 -5041 140167 -5007
rect 142003 -5041 142015 -5007
rect 143851 -5041 143863 -5007
rect 145699 -5041 145711 -5007
rect 147547 -5041 147559 -5007
rect 149395 -5041 149407 -5007
rect 151243 -5041 151255 -5007
rect 153091 -5041 153103 -5007
rect 154939 -5041 154951 -5007
rect 156787 -5041 156799 -5007
rect 158635 -5041 158647 -5007
rect 160483 -5041 160495 -5007
rect 162331 -5041 162343 -5007
rect 164179 -5041 164191 -5007
rect 166027 -5041 166039 -5007
rect 167875 -5041 167887 -5007
rect 169723 -5041 169735 -5007
rect 171571 -5041 171583 -5007
rect 173419 -5041 173431 -5007
rect 175267 -5041 175279 -5007
rect 177115 -5041 177127 -5007
rect 178963 -5041 178975 -5007
rect 3403 -5047 3461 -5041
rect 5251 -5047 5309 -5041
rect 7099 -5047 7157 -5041
rect 8947 -5047 9005 -5041
rect 10795 -5047 10853 -5041
rect 12643 -5047 12701 -5041
rect 14491 -5047 14549 -5041
rect 16339 -5047 16397 -5041
rect 18187 -5047 18245 -5041
rect 20035 -5047 20093 -5041
rect 21883 -5047 21941 -5041
rect 23731 -5047 23789 -5041
rect 25579 -5047 25637 -5041
rect 27427 -5047 27485 -5041
rect 29275 -5047 29333 -5041
rect 31123 -5047 31181 -5041
rect 32971 -5047 33029 -5041
rect 34819 -5047 34877 -5041
rect 36667 -5047 36725 -5041
rect 38515 -5047 38573 -5041
rect 40363 -5047 40421 -5041
rect 42211 -5047 42269 -5041
rect 44059 -5047 44117 -5041
rect 45907 -5047 45965 -5041
rect 47755 -5047 47813 -5041
rect 49603 -5047 49661 -5041
rect 51451 -5047 51509 -5041
rect 53299 -5047 53357 -5041
rect 55147 -5047 55205 -5041
rect 56995 -5047 57053 -5041
rect 58843 -5047 58901 -5041
rect 60691 -5047 60749 -5041
rect 62539 -5047 62597 -5041
rect 64387 -5047 64445 -5041
rect 66235 -5047 66293 -5041
rect 68083 -5047 68141 -5041
rect 69931 -5047 69989 -5041
rect 71779 -5047 71837 -5041
rect 73627 -5047 73685 -5041
rect 75475 -5047 75533 -5041
rect 77323 -5047 77381 -5041
rect 79171 -5047 79229 -5041
rect 81019 -5047 81077 -5041
rect 82867 -5047 82925 -5041
rect 84715 -5047 84773 -5041
rect 86563 -5047 86621 -5041
rect 88411 -5047 88469 -5041
rect 90259 -5047 90317 -5041
rect 92107 -5047 92165 -5041
rect 93955 -5047 94013 -5041
rect 95803 -5047 95861 -5041
rect 97651 -5047 97709 -5041
rect 99499 -5047 99557 -5041
rect 101347 -5047 101405 -5041
rect 103195 -5047 103253 -5041
rect 105043 -5047 105101 -5041
rect 106891 -5047 106949 -5041
rect 108739 -5047 108797 -5041
rect 110587 -5047 110645 -5041
rect 112435 -5047 112493 -5041
rect 114283 -5047 114341 -5041
rect 116131 -5047 116189 -5041
rect 117979 -5047 118037 -5041
rect 119827 -5047 119885 -5041
rect 121675 -5047 121733 -5041
rect 123523 -5047 123581 -5041
rect 125371 -5047 125429 -5041
rect 127219 -5047 127277 -5041
rect 129067 -5047 129125 -5041
rect 130915 -5047 130973 -5041
rect 132763 -5047 132821 -5041
rect 134611 -5047 134669 -5041
rect 136459 -5047 136517 -5041
rect 138307 -5047 138365 -5041
rect 140155 -5047 140213 -5041
rect 142003 -5047 142061 -5041
rect 143851 -5047 143909 -5041
rect 145699 -5047 145757 -5041
rect 147547 -5047 147605 -5041
rect 149395 -5047 149453 -5041
rect 151243 -5047 151301 -5041
rect 153091 -5047 153149 -5041
rect 154939 -5047 154997 -5041
rect 156787 -5047 156845 -5041
rect 158635 -5047 158693 -5041
rect 160483 -5047 160541 -5041
rect 162331 -5047 162389 -5041
rect 164179 -5047 164237 -5041
rect 166027 -5047 166085 -5041
rect 167875 -5047 167933 -5041
rect 169723 -5047 169781 -5041
rect 171571 -5047 171629 -5041
rect 173419 -5047 173477 -5041
rect 175267 -5047 175325 -5041
rect 177115 -5047 177173 -5041
rect 178963 -5047 179021 -5041
rect 413 -5229 659 -5196
rect 1555 -5201 1613 -5195
rect 3403 -5201 3461 -5195
rect 5251 -5201 5309 -5195
rect 7099 -5201 7157 -5195
rect 8947 -5201 9005 -5195
rect 10795 -5201 10853 -5195
rect 12643 -5201 12701 -5195
rect 14491 -5201 14549 -5195
rect 16339 -5201 16397 -5195
rect 18187 -5201 18245 -5195
rect 20035 -5201 20093 -5195
rect 21883 -5201 21941 -5195
rect 23731 -5201 23789 -5195
rect 25579 -5201 25637 -5195
rect 27427 -5201 27485 -5195
rect 29275 -5201 29333 -5195
rect 31123 -5201 31181 -5195
rect 32971 -5201 33029 -5195
rect 34819 -5201 34877 -5195
rect 36667 -5201 36725 -5195
rect 38515 -5201 38573 -5195
rect 40363 -5201 40421 -5195
rect 42211 -5201 42269 -5195
rect 44059 -5201 44117 -5195
rect 45907 -5201 45965 -5195
rect 47755 -5201 47813 -5195
rect 49603 -5201 49661 -5195
rect 51451 -5201 51509 -5195
rect 53299 -5201 53357 -5195
rect 55147 -5201 55205 -5195
rect 56995 -5201 57053 -5195
rect 58843 -5201 58901 -5195
rect 60691 -5201 60749 -5195
rect 62539 -5201 62597 -5195
rect 64387 -5201 64445 -5195
rect 66235 -5201 66293 -5195
rect 68083 -5201 68141 -5195
rect 69931 -5201 69989 -5195
rect 71779 -5201 71837 -5195
rect 73627 -5201 73685 -5195
rect 75475 -5201 75533 -5195
rect 77323 -5201 77381 -5195
rect 79171 -5201 79229 -5195
rect 81019 -5201 81077 -5195
rect 82867 -5201 82925 -5195
rect 84715 -5201 84773 -5195
rect 86563 -5201 86621 -5195
rect 88411 -5201 88469 -5195
rect 90259 -5201 90317 -5195
rect 92107 -5201 92165 -5195
rect 93955 -5201 94013 -5195
rect 95803 -5201 95861 -5195
rect 97651 -5201 97709 -5195
rect 99499 -5201 99557 -5195
rect 101347 -5201 101405 -5195
rect 103195 -5201 103253 -5195
rect 105043 -5201 105101 -5195
rect 106891 -5201 106949 -5195
rect 108739 -5201 108797 -5195
rect 110587 -5201 110645 -5195
rect 112435 -5201 112493 -5195
rect 114283 -5201 114341 -5195
rect 116131 -5201 116189 -5195
rect 117979 -5201 118037 -5195
rect 119827 -5201 119885 -5195
rect 121675 -5201 121733 -5195
rect 123523 -5201 123581 -5195
rect 125371 -5201 125429 -5195
rect 127219 -5201 127277 -5195
rect 129067 -5201 129125 -5195
rect 130915 -5201 130973 -5195
rect 132763 -5201 132821 -5195
rect 134611 -5201 134669 -5195
rect 136459 -5201 136517 -5195
rect 138307 -5201 138365 -5195
rect 140155 -5201 140213 -5195
rect 142003 -5201 142061 -5195
rect 143851 -5201 143909 -5195
rect 145699 -5201 145757 -5195
rect 147547 -5201 147605 -5195
rect 149395 -5201 149453 -5195
rect 151243 -5201 151301 -5195
rect 153091 -5201 153149 -5195
rect 154939 -5201 154997 -5195
rect 156787 -5201 156845 -5195
rect 158635 -5201 158693 -5195
rect 160483 -5201 160541 -5195
rect 162331 -5201 162389 -5195
rect 164179 -5201 164237 -5195
rect 166027 -5201 166085 -5195
rect 167875 -5201 167933 -5195
rect 169723 -5201 169781 -5195
rect 171571 -5201 171629 -5195
rect 173419 -5201 173477 -5195
rect 175267 -5201 175325 -5195
rect 177115 -5201 177173 -5195
rect 178963 -5201 179021 -5195
rect 396 -5232 659 -5229
rect 976 -5232 1028 -5231
rect 296 -5247 307 -5236
rect 222 -5257 307 -5247
rect 80 -5263 307 -5257
rect 396 -5263 896 -5232
rect 80 -5266 896 -5263
rect 80 -5297 659 -5266
rect 958 -5267 1028 -5232
rect 80 -5345 307 -5297
rect 396 -5318 659 -5297
rect 833 -5300 880 -5287
rect 665 -5318 676 -5307
rect 396 -5334 676 -5318
rect 765 -5328 880 -5300
rect 976 -5328 1046 -5267
rect 1108 -5301 1267 -5267
rect 1327 -5301 1363 -5284
rect 765 -5334 1046 -5328
rect 396 -5345 1046 -5334
rect 1328 -5302 1363 -5301
rect 1373 -5302 1399 -5231
rect 1328 -5338 1399 -5302
rect 1409 -5284 1417 -5213
rect 1555 -5235 1567 -5201
rect 3403 -5235 3415 -5201
rect 5251 -5235 5263 -5201
rect 7099 -5235 7111 -5201
rect 8947 -5235 8959 -5201
rect 10795 -5235 10807 -5201
rect 12643 -5235 12655 -5201
rect 14491 -5235 14503 -5201
rect 16339 -5235 16351 -5201
rect 18187 -5235 18199 -5201
rect 20035 -5235 20047 -5201
rect 21883 -5235 21895 -5201
rect 23731 -5235 23743 -5201
rect 25579 -5235 25591 -5201
rect 27427 -5235 27439 -5201
rect 29275 -5235 29287 -5201
rect 31123 -5235 31135 -5201
rect 32971 -5235 32983 -5201
rect 34819 -5235 34831 -5201
rect 36667 -5235 36679 -5201
rect 38515 -5235 38527 -5201
rect 40363 -5235 40375 -5201
rect 42211 -5235 42223 -5201
rect 44059 -5235 44071 -5201
rect 45907 -5235 45919 -5201
rect 47755 -5235 47767 -5201
rect 49603 -5235 49615 -5201
rect 51451 -5235 51463 -5201
rect 53299 -5235 53311 -5201
rect 55147 -5235 55159 -5201
rect 56995 -5235 57007 -5201
rect 58843 -5235 58855 -5201
rect 60691 -5235 60703 -5201
rect 62539 -5235 62551 -5201
rect 64387 -5235 64399 -5201
rect 66235 -5235 66247 -5201
rect 68083 -5235 68095 -5201
rect 69931 -5235 69943 -5201
rect 71779 -5235 71791 -5201
rect 73627 -5235 73639 -5201
rect 75475 -5235 75487 -5201
rect 77323 -5235 77335 -5201
rect 79171 -5235 79183 -5201
rect 81019 -5235 81031 -5201
rect 82867 -5235 82879 -5201
rect 84715 -5235 84727 -5201
rect 86563 -5235 86575 -5201
rect 88411 -5235 88423 -5201
rect 90259 -5235 90271 -5201
rect 92107 -5235 92119 -5201
rect 93955 -5235 93967 -5201
rect 95803 -5235 95815 -5201
rect 97651 -5235 97663 -5201
rect 99499 -5235 99511 -5201
rect 101347 -5235 101359 -5201
rect 103195 -5235 103207 -5201
rect 105043 -5235 105055 -5201
rect 106891 -5235 106903 -5201
rect 108739 -5235 108751 -5201
rect 110587 -5235 110599 -5201
rect 112435 -5235 112447 -5201
rect 114283 -5235 114295 -5201
rect 116131 -5235 116143 -5201
rect 117979 -5235 117991 -5201
rect 119827 -5235 119839 -5201
rect 121675 -5235 121687 -5201
rect 123523 -5235 123535 -5201
rect 125371 -5235 125383 -5201
rect 127219 -5235 127231 -5201
rect 129067 -5235 129079 -5201
rect 130915 -5235 130927 -5201
rect 132763 -5235 132775 -5201
rect 134611 -5235 134623 -5201
rect 136459 -5235 136471 -5201
rect 138307 -5235 138319 -5201
rect 140155 -5235 140167 -5201
rect 142003 -5235 142015 -5201
rect 143851 -5235 143863 -5201
rect 145699 -5235 145711 -5201
rect 147547 -5235 147559 -5201
rect 149395 -5235 149407 -5201
rect 151243 -5235 151255 -5201
rect 153091 -5235 153103 -5201
rect 154939 -5235 154951 -5201
rect 156787 -5235 156799 -5201
rect 158635 -5235 158647 -5201
rect 160483 -5235 160495 -5201
rect 162331 -5235 162343 -5201
rect 164179 -5235 164191 -5201
rect 166027 -5235 166039 -5201
rect 167875 -5235 167887 -5201
rect 169723 -5235 169735 -5201
rect 171571 -5235 171583 -5201
rect 173419 -5235 173431 -5201
rect 175267 -5235 175279 -5201
rect 177115 -5235 177127 -5201
rect 178963 -5235 178975 -5201
rect 1555 -5241 1613 -5235
rect 3403 -5241 3461 -5235
rect 5251 -5241 5309 -5235
rect 7099 -5241 7157 -5235
rect 8947 -5241 9005 -5235
rect 10795 -5241 10853 -5235
rect 12643 -5241 12701 -5235
rect 14491 -5241 14549 -5235
rect 16339 -5241 16397 -5235
rect 18187 -5241 18245 -5235
rect 20035 -5241 20093 -5235
rect 21883 -5241 21941 -5235
rect 23731 -5241 23789 -5235
rect 25579 -5241 25637 -5235
rect 27427 -5241 27485 -5235
rect 29275 -5241 29333 -5235
rect 31123 -5241 31181 -5235
rect 32971 -5241 33029 -5235
rect 34819 -5241 34877 -5235
rect 36667 -5241 36725 -5235
rect 38515 -5241 38573 -5235
rect 40363 -5241 40421 -5235
rect 42211 -5241 42269 -5235
rect 44059 -5241 44117 -5235
rect 45907 -5241 45965 -5235
rect 47755 -5241 47813 -5235
rect 49603 -5241 49661 -5235
rect 51451 -5241 51509 -5235
rect 53299 -5241 53357 -5235
rect 55147 -5241 55205 -5235
rect 56995 -5241 57053 -5235
rect 58843 -5241 58901 -5235
rect 60691 -5241 60749 -5235
rect 62539 -5241 62597 -5235
rect 64387 -5241 64445 -5235
rect 66235 -5241 66293 -5235
rect 68083 -5241 68141 -5235
rect 69931 -5241 69989 -5235
rect 71779 -5241 71837 -5235
rect 73627 -5241 73685 -5235
rect 75475 -5241 75533 -5235
rect 77323 -5241 77381 -5235
rect 79171 -5241 79229 -5235
rect 81019 -5241 81077 -5235
rect 82867 -5241 82925 -5235
rect 84715 -5241 84773 -5235
rect 86563 -5241 86621 -5235
rect 88411 -5241 88469 -5235
rect 90259 -5241 90317 -5235
rect 92107 -5241 92165 -5235
rect 93955 -5241 94013 -5235
rect 95803 -5241 95861 -5235
rect 97651 -5241 97709 -5235
rect 99499 -5241 99557 -5235
rect 101347 -5241 101405 -5235
rect 103195 -5241 103253 -5235
rect 105043 -5241 105101 -5235
rect 106891 -5241 106949 -5235
rect 108739 -5241 108797 -5235
rect 110587 -5241 110645 -5235
rect 112435 -5241 112493 -5235
rect 114283 -5241 114341 -5235
rect 116131 -5241 116189 -5235
rect 117979 -5241 118037 -5235
rect 119827 -5241 119885 -5235
rect 121675 -5241 121733 -5235
rect 123523 -5241 123581 -5235
rect 125371 -5241 125429 -5235
rect 127219 -5241 127277 -5235
rect 129067 -5241 129125 -5235
rect 130915 -5241 130973 -5235
rect 132763 -5241 132821 -5235
rect 134611 -5241 134669 -5235
rect 136459 -5241 136517 -5235
rect 138307 -5241 138365 -5235
rect 140155 -5241 140213 -5235
rect 142003 -5241 142061 -5235
rect 143851 -5241 143909 -5235
rect 145699 -5241 145757 -5235
rect 147547 -5241 147605 -5235
rect 149395 -5241 149453 -5235
rect 151243 -5241 151301 -5235
rect 153091 -5241 153149 -5235
rect 154939 -5241 154997 -5235
rect 156787 -5241 156845 -5235
rect 158635 -5241 158693 -5235
rect 160483 -5241 160541 -5235
rect 162331 -5241 162389 -5235
rect 164179 -5241 164237 -5235
rect 166027 -5241 166085 -5235
rect 167875 -5241 167933 -5235
rect 169723 -5241 169781 -5235
rect 171571 -5241 171629 -5235
rect 173419 -5241 173477 -5235
rect 175267 -5241 175325 -5235
rect 177115 -5241 177173 -5235
rect 178963 -5241 179021 -5235
rect 1409 -5303 1443 -5284
rect 1725 -5303 1759 -5284
rect 1409 -5337 1759 -5303
rect 1716 -5338 1795 -5337
rect 80 -5363 1046 -5345
rect 1345 -5363 1795 -5338
rect 80 -5368 1047 -5363
rect 80 -5389 676 -5368
rect 79 -5407 676 -5389
rect 765 -5407 1047 -5368
rect 79 -5422 1047 -5407
rect 1158 -5369 1217 -5363
rect 1158 -5403 1205 -5369
rect 1328 -5371 1795 -5363
rect 1328 -5372 1417 -5371
rect 1477 -5372 1636 -5371
rect 1158 -5409 1217 -5403
rect 79 -5423 333 -5422
rect 80 -5481 333 -5423
rect 396 -5481 1047 -5422
rect 80 -5484 1047 -5481
rect 80 -5521 676 -5484
rect 125 -5525 213 -5521
rect 125 -5541 191 -5525
rect 222 -5531 676 -5521
rect 298 -5534 676 -5531
rect 765 -5534 1047 -5484
rect 1126 -5528 1161 -5462
rect 1214 -5528 1249 -5462
rect 143 -5550 173 -5541
rect 298 -5550 1047 -5534
rect 143 -5572 253 -5550
rect 85 -5583 253 -5572
rect 299 -5568 1047 -5550
rect 299 -5583 702 -5568
rect 85 -5584 702 -5583
rect 85 -5617 659 -5584
rect 691 -5595 702 -5584
rect 765 -5574 1047 -5568
rect 765 -5584 850 -5574
rect 765 -5595 776 -5584
rect 299 -5636 659 -5617
rect 976 -5627 1047 -5574
rect 1170 -5621 1205 -5587
rect 1328 -5627 1416 -5372
rect 1698 -5373 1795 -5371
rect 1716 -5434 1786 -5373
rect 1848 -5389 2007 -5373
rect 1848 -5390 2085 -5389
rect 1848 -5407 2147 -5390
rect 1527 -5440 1586 -5434
rect 1527 -5474 1574 -5440
rect 1697 -5469 1786 -5434
rect 1527 -5480 1586 -5474
rect 1495 -5590 1530 -5524
rect 1583 -5590 1618 -5524
rect 299 -5653 896 -5636
rect 299 -5839 386 -5653
rect 494 -5659 896 -5653
rect 483 -5670 896 -5659
rect 976 -5670 1046 -5627
rect 498 -5686 510 -5670
rect 498 -5692 556 -5686
rect 316 -5935 386 -5839
rect 498 -5852 556 -5846
rect 498 -5886 510 -5852
rect 498 -5892 556 -5886
rect 668 -5892 702 -5670
rect 976 -5706 1028 -5670
rect 1108 -5723 1267 -5689
rect 1345 -5723 1416 -5627
rect 1527 -5640 1586 -5634
rect 1527 -5674 1574 -5640
rect 1527 -5680 1586 -5674
rect 1697 -5680 1787 -5469
rect 1345 -5759 1399 -5723
rect 1716 -5733 1787 -5680
rect 1831 -5485 1841 -5407
rect 1927 -5408 2147 -5407
rect 1927 -5423 2217 -5408
rect 1860 -5485 1865 -5441
rect 2068 -5444 2217 -5423
rect 2456 -5444 2508 -5443
rect 1931 -5475 1961 -5459
rect 2085 -5469 2376 -5444
rect 1477 -5776 1636 -5742
rect 1716 -5776 1786 -5733
rect 1716 -5812 1768 -5776
rect 1831 -5795 1865 -5485
rect 1894 -5509 1899 -5475
rect 1910 -5509 1961 -5475
rect 1973 -5518 2003 -5475
rect 2068 -5478 2376 -5469
rect 1973 -5525 2023 -5518
rect 2034 -5525 2039 -5491
rect 1973 -5528 1985 -5525
rect 1973 -5531 2023 -5528
rect 1973 -5541 1985 -5531
rect 1975 -5552 1991 -5546
rect 1866 -5568 1899 -5552
rect 1954 -5556 1991 -5552
rect 2068 -5550 2217 -5478
rect 2438 -5479 2508 -5444
rect 2456 -5514 2526 -5479
rect 2588 -5496 2750 -5479
rect 2530 -5513 2750 -5496
rect 2807 -5513 2846 -5496
rect 2808 -5514 2846 -5513
rect 3995 -5514 4029 -5496
rect 5843 -5514 5877 -5496
rect 7691 -5514 7725 -5496
rect 9539 -5514 9573 -5496
rect 11387 -5514 11421 -5496
rect 13235 -5514 13269 -5496
rect 15083 -5514 15117 -5496
rect 16931 -5514 16965 -5496
rect 18779 -5514 18813 -5496
rect 20627 -5514 20661 -5496
rect 22475 -5514 22509 -5496
rect 24323 -5514 24357 -5496
rect 26171 -5514 26205 -5496
rect 28019 -5514 28053 -5496
rect 29867 -5514 29901 -5496
rect 31715 -5514 31749 -5496
rect 33563 -5514 33597 -5496
rect 35411 -5514 35445 -5496
rect 37259 -5514 37293 -5496
rect 39107 -5514 39141 -5496
rect 40955 -5514 40989 -5496
rect 42803 -5514 42837 -5496
rect 44651 -5514 44685 -5496
rect 46499 -5514 46533 -5496
rect 48347 -5514 48381 -5496
rect 50195 -5514 50229 -5496
rect 52043 -5514 52077 -5496
rect 53891 -5514 53925 -5496
rect 55739 -5514 55773 -5496
rect 57587 -5514 57621 -5496
rect 59435 -5514 59469 -5496
rect 61283 -5514 61317 -5496
rect 63131 -5514 63165 -5496
rect 64979 -5514 65013 -5496
rect 66827 -5514 66861 -5496
rect 68675 -5514 68709 -5496
rect 70523 -5514 70557 -5496
rect 72371 -5514 72405 -5496
rect 74219 -5514 74253 -5496
rect 76067 -5514 76101 -5496
rect 77915 -5514 77949 -5496
rect 79763 -5514 79797 -5496
rect 81611 -5514 81645 -5496
rect 83459 -5514 83493 -5496
rect 85307 -5514 85341 -5496
rect 87155 -5514 87189 -5496
rect 89003 -5514 89037 -5496
rect 90851 -5514 90885 -5496
rect 92699 -5514 92733 -5496
rect 94547 -5514 94581 -5496
rect 96395 -5514 96429 -5496
rect 98243 -5514 98277 -5496
rect 100091 -5514 100125 -5496
rect 101939 -5514 101973 -5496
rect 103787 -5514 103821 -5496
rect 105635 -5514 105669 -5496
rect 107483 -5514 107517 -5496
rect 109331 -5514 109365 -5496
rect 111179 -5514 111213 -5496
rect 113027 -5514 113061 -5496
rect 114875 -5514 114909 -5496
rect 116723 -5514 116757 -5496
rect 118571 -5514 118605 -5496
rect 120419 -5514 120453 -5496
rect 122267 -5514 122301 -5496
rect 124115 -5514 124149 -5496
rect 125963 -5514 125997 -5496
rect 127811 -5514 127845 -5496
rect 129659 -5514 129693 -5496
rect 131507 -5514 131541 -5496
rect 133355 -5514 133389 -5496
rect 135203 -5514 135237 -5496
rect 137051 -5514 137085 -5496
rect 138899 -5514 138933 -5496
rect 140747 -5514 140781 -5496
rect 142595 -5514 142629 -5496
rect 144443 -5514 144477 -5496
rect 146291 -5514 146325 -5496
rect 148139 -5514 148173 -5496
rect 149987 -5514 150021 -5496
rect 151835 -5514 151869 -5496
rect 153683 -5514 153717 -5496
rect 155531 -5514 155565 -5496
rect 157379 -5514 157413 -5496
rect 159227 -5514 159261 -5496
rect 161075 -5514 161109 -5496
rect 162923 -5514 162957 -5496
rect 164771 -5514 164805 -5496
rect 166619 -5514 166653 -5496
rect 168467 -5514 168501 -5496
rect 170315 -5514 170349 -5496
rect 172163 -5514 172197 -5496
rect 174011 -5514 174045 -5496
rect 175859 -5514 175893 -5496
rect 177707 -5514 177741 -5496
rect 179501 -5513 179536 -5496
rect 179502 -5514 179536 -5513
rect 179924 -5513 179959 -5496
rect 180239 -5513 180274 -5496
rect 179924 -5514 179958 -5513
rect 2456 -5540 2586 -5514
rect 2267 -5546 2326 -5540
rect 2267 -5550 2314 -5546
rect 2437 -5550 2586 -5540
rect 2808 -5550 2882 -5514
rect 3995 -5550 4065 -5514
rect 5843 -5550 5913 -5514
rect 7691 -5550 7761 -5514
rect 9539 -5550 9609 -5514
rect 11387 -5550 11457 -5514
rect 13235 -5550 13305 -5514
rect 15083 -5550 15153 -5514
rect 16931 -5550 17001 -5514
rect 18779 -5550 18849 -5514
rect 20627 -5550 20697 -5514
rect 22475 -5550 22545 -5514
rect 24323 -5550 24393 -5514
rect 26171 -5550 26241 -5514
rect 28019 -5550 28089 -5514
rect 29867 -5550 29937 -5514
rect 31715 -5550 31785 -5514
rect 33563 -5550 33633 -5514
rect 35411 -5550 35481 -5514
rect 37259 -5550 37329 -5514
rect 39107 -5550 39177 -5514
rect 40955 -5550 41025 -5514
rect 42803 -5550 42873 -5514
rect 44651 -5550 44721 -5514
rect 46499 -5550 46569 -5514
rect 48347 -5550 48417 -5514
rect 50195 -5550 50265 -5514
rect 52043 -5550 52113 -5514
rect 53891 -5550 53961 -5514
rect 55739 -5550 55809 -5514
rect 57587 -5550 57657 -5514
rect 59435 -5550 59505 -5514
rect 61283 -5550 61353 -5514
rect 63131 -5550 63201 -5514
rect 64979 -5550 65049 -5514
rect 66827 -5550 66897 -5514
rect 68675 -5550 68745 -5514
rect 70523 -5550 70593 -5514
rect 72371 -5550 72441 -5514
rect 74219 -5550 74289 -5514
rect 76067 -5550 76137 -5514
rect 77915 -5550 77985 -5514
rect 79763 -5550 79833 -5514
rect 81611 -5550 81681 -5514
rect 83459 -5550 83529 -5514
rect 85307 -5550 85377 -5514
rect 87155 -5550 87225 -5514
rect 89003 -5550 89073 -5514
rect 90851 -5550 90921 -5514
rect 92699 -5550 92769 -5514
rect 94547 -5550 94617 -5514
rect 96395 -5550 96465 -5514
rect 98243 -5550 98313 -5514
rect 100091 -5550 100161 -5514
rect 101939 -5550 102009 -5514
rect 103787 -5550 103857 -5514
rect 105635 -5550 105705 -5514
rect 107483 -5550 107553 -5514
rect 109331 -5550 109401 -5514
rect 111179 -5550 111249 -5514
rect 113027 -5550 113097 -5514
rect 114875 -5550 114945 -5514
rect 116723 -5550 116793 -5514
rect 118571 -5550 118641 -5514
rect 120419 -5550 120489 -5514
rect 122267 -5550 122337 -5514
rect 124115 -5550 124185 -5514
rect 125963 -5550 126033 -5514
rect 127811 -5550 127881 -5514
rect 129659 -5550 129729 -5514
rect 131507 -5550 131577 -5514
rect 133355 -5550 133425 -5514
rect 135203 -5550 135273 -5514
rect 137051 -5550 137121 -5514
rect 138899 -5550 138969 -5514
rect 140747 -5550 140817 -5514
rect 142595 -5550 142665 -5514
rect 144443 -5550 144513 -5514
rect 146291 -5550 146361 -5514
rect 148139 -5550 148209 -5514
rect 149987 -5550 150057 -5514
rect 151835 -5550 151905 -5514
rect 153683 -5550 153753 -5514
rect 155531 -5550 155601 -5514
rect 157379 -5550 157449 -5514
rect 159227 -5550 159297 -5514
rect 161075 -5550 161145 -5514
rect 162923 -5550 162993 -5514
rect 164771 -5550 164841 -5514
rect 166619 -5550 166689 -5514
rect 168467 -5550 168537 -5514
rect 170315 -5550 170385 -5514
rect 172163 -5550 172233 -5514
rect 174011 -5550 174081 -5514
rect 175859 -5550 175929 -5514
rect 177707 -5550 177777 -5514
rect 179502 -5550 179572 -5514
rect 1949 -5559 2001 -5556
rect 1975 -5568 2001 -5559
rect 2068 -5564 2235 -5550
rect 2252 -5561 2586 -5550
rect 2263 -5564 2586 -5561
rect 1866 -5634 1901 -5568
rect 1954 -5572 2001 -5568
rect 1934 -5584 1943 -5573
rect 1954 -5584 1989 -5572
rect 1945 -5634 1989 -5584
rect 1991 -5634 2000 -5572
rect 1866 -5650 1899 -5634
rect 1945 -5646 1979 -5634
rect 1933 -5672 1979 -5646
rect 1933 -5677 1943 -5672
rect 1945 -5677 1979 -5672
rect 1933 -5693 1979 -5677
rect 1894 -5727 1899 -5693
rect 1910 -5727 1979 -5693
rect 1933 -5740 1979 -5727
rect 1933 -5741 1961 -5740
rect 2034 -5741 2067 -5568
rect 2068 -5584 2586 -5564
rect 2825 -5575 2900 -5550
rect 2068 -5618 2234 -5584
rect 2267 -5586 2326 -5584
rect 2235 -5618 2270 -5614
rect 2323 -5618 2358 -5614
rect 2068 -5630 2268 -5618
rect 2355 -5630 2370 -5621
rect 2068 -5696 2270 -5630
rect 2323 -5670 2370 -5630
rect 2068 -5708 2268 -5696
rect 2312 -5708 2370 -5670
rect 2403 -5686 2408 -5652
rect 2068 -5741 2234 -5708
rect 2235 -5712 2268 -5708
rect 2323 -5712 2358 -5708
rect 2314 -5724 2348 -5720
rect 1933 -5752 1973 -5741
rect 2034 -5752 2234 -5741
rect 2302 -5736 2354 -5724
rect 2302 -5746 2348 -5736
rect 2034 -5756 2067 -5752
rect 1955 -5795 2007 -5765
rect 2068 -5790 2234 -5752
rect 2263 -5780 2268 -5746
rect 2279 -5780 2330 -5746
rect 1831 -5829 2061 -5795
rect 1831 -5839 1865 -5829
rect 2085 -5848 2234 -5790
rect 2302 -5794 2330 -5780
rect 2403 -5794 2436 -5720
rect 2437 -5794 2586 -5584
rect 2638 -5581 2700 -5575
rect 2638 -5615 2688 -5581
rect 2808 -5584 2900 -5575
rect 2957 -5584 3119 -5550
rect 4012 -5584 4083 -5550
rect 5860 -5584 5931 -5550
rect 7708 -5584 7779 -5550
rect 9556 -5584 9627 -5550
rect 11404 -5584 11475 -5550
rect 13252 -5584 13323 -5550
rect 15100 -5584 15171 -5550
rect 16948 -5584 17019 -5550
rect 18796 -5584 18867 -5550
rect 20644 -5584 20715 -5550
rect 22492 -5584 22563 -5550
rect 24340 -5584 24411 -5550
rect 26188 -5584 26259 -5550
rect 28036 -5584 28107 -5550
rect 29884 -5584 29955 -5550
rect 31732 -5584 31803 -5550
rect 33580 -5584 33651 -5550
rect 35428 -5584 35499 -5550
rect 37276 -5584 37347 -5550
rect 39124 -5584 39195 -5550
rect 40972 -5584 41043 -5550
rect 42820 -5584 42891 -5550
rect 44668 -5584 44739 -5550
rect 46516 -5584 46587 -5550
rect 48364 -5584 48435 -5550
rect 50212 -5584 50283 -5550
rect 52060 -5584 52131 -5550
rect 53908 -5584 53979 -5550
rect 55756 -5584 55827 -5550
rect 57604 -5584 57675 -5550
rect 59452 -5584 59523 -5550
rect 61300 -5584 61371 -5550
rect 63148 -5584 63219 -5550
rect 64996 -5584 65067 -5550
rect 66844 -5584 66915 -5550
rect 68692 -5584 68763 -5550
rect 70540 -5584 70611 -5550
rect 72388 -5584 72459 -5550
rect 74236 -5584 74307 -5550
rect 76084 -5584 76155 -5550
rect 77932 -5584 78003 -5550
rect 79780 -5584 79851 -5550
rect 81628 -5584 81699 -5550
rect 83476 -5584 83547 -5550
rect 85324 -5584 85395 -5550
rect 87172 -5584 87243 -5550
rect 89020 -5584 89091 -5550
rect 90868 -5584 90939 -5550
rect 92716 -5584 92787 -5550
rect 94564 -5584 94635 -5550
rect 96412 -5584 96483 -5550
rect 98260 -5584 98331 -5550
rect 100108 -5584 100179 -5550
rect 101956 -5584 102027 -5550
rect 103804 -5584 103875 -5550
rect 105652 -5584 105723 -5550
rect 107500 -5584 107571 -5550
rect 109348 -5584 109419 -5550
rect 111196 -5584 111267 -5550
rect 113044 -5584 113115 -5550
rect 114892 -5584 114963 -5550
rect 116740 -5584 116811 -5550
rect 118588 -5584 118659 -5550
rect 120436 -5584 120507 -5550
rect 122284 -5584 122355 -5550
rect 124132 -5584 124203 -5550
rect 125980 -5584 126051 -5550
rect 127828 -5584 127899 -5550
rect 129676 -5584 129747 -5550
rect 131524 -5584 131595 -5550
rect 133372 -5584 133443 -5550
rect 135220 -5584 135291 -5550
rect 137068 -5584 137139 -5550
rect 138916 -5584 138987 -5550
rect 140764 -5584 140835 -5550
rect 142612 -5584 142683 -5550
rect 144460 -5584 144531 -5550
rect 146308 -5584 146379 -5550
rect 148156 -5584 148227 -5550
rect 150004 -5584 150075 -5550
rect 151852 -5584 151923 -5550
rect 153700 -5584 153771 -5550
rect 155548 -5584 155619 -5550
rect 157396 -5584 157467 -5550
rect 159244 -5584 159315 -5550
rect 161092 -5584 161163 -5550
rect 162940 -5584 163011 -5550
rect 164788 -5584 164859 -5550
rect 166636 -5584 166707 -5550
rect 168484 -5584 168555 -5550
rect 170332 -5584 170403 -5550
rect 172180 -5584 172251 -5550
rect 174028 -5584 174099 -5550
rect 175876 -5584 175947 -5550
rect 177724 -5584 177795 -5550
rect 179332 -5581 179390 -5575
rect 2638 -5621 2700 -5615
rect 2594 -5752 2604 -5662
rect 2606 -5740 2644 -5674
rect 2652 -5740 2655 -5663
rect 2683 -5674 2686 -5663
rect 2694 -5740 2732 -5674
rect 2302 -5814 2342 -5794
rect 2403 -5814 2586 -5794
rect 2314 -5818 2348 -5814
rect 2402 -5818 2436 -5814
rect 2324 -5846 2376 -5818
rect 2324 -5848 2404 -5846
rect 2437 -5848 2586 -5814
rect 2650 -5833 2688 -5799
rect 2808 -5839 2899 -5584
rect 3007 -5652 3069 -5646
rect 3007 -5686 3057 -5652
rect 3007 -5692 3069 -5686
rect 2975 -5802 3013 -5736
rect 3021 -5802 3024 -5725
rect 3052 -5736 3055 -5725
rect 3063 -5802 3101 -5736
rect 2085 -5852 2586 -5848
rect 2085 -5882 2439 -5852
rect 2085 -5918 2234 -5882
rect 2346 -5886 2358 -5882
rect 2346 -5892 2404 -5886
rect 2164 -5935 2234 -5918
rect 316 -5971 369 -5935
rect 2164 -5971 2217 -5935
rect 2456 -5971 2586 -5852
rect 2588 -5935 2750 -5901
rect 2825 -5935 2899 -5839
rect 3007 -5852 3069 -5846
rect 3007 -5886 3057 -5852
rect 3007 -5892 3069 -5886
rect 3177 -5892 3215 -5646
rect 4012 -5935 4082 -5584
rect 4194 -5652 4252 -5646
rect 4194 -5686 4206 -5652
rect 4194 -5692 4252 -5686
rect 4194 -5852 4252 -5846
rect 4194 -5886 4206 -5852
rect 4194 -5892 4252 -5886
rect 5860 -5935 5930 -5584
rect 6042 -5652 6100 -5646
rect 6042 -5686 6054 -5652
rect 6042 -5692 6100 -5686
rect 6042 -5852 6100 -5846
rect 6042 -5886 6054 -5852
rect 6042 -5892 6100 -5886
rect 7708 -5935 7778 -5584
rect 7890 -5652 7948 -5646
rect 7890 -5686 7902 -5652
rect 7890 -5692 7948 -5686
rect 7890 -5852 7948 -5846
rect 7890 -5886 7902 -5852
rect 7890 -5892 7948 -5886
rect 9556 -5935 9626 -5584
rect 9738 -5652 9796 -5646
rect 9738 -5686 9750 -5652
rect 9738 -5692 9796 -5686
rect 9738 -5852 9796 -5846
rect 9738 -5886 9750 -5852
rect 9738 -5892 9796 -5886
rect 11404 -5935 11474 -5584
rect 11586 -5652 11644 -5646
rect 11586 -5686 11598 -5652
rect 11586 -5692 11644 -5686
rect 11586 -5852 11644 -5846
rect 11586 -5886 11598 -5852
rect 11586 -5892 11644 -5886
rect 13252 -5935 13322 -5584
rect 13434 -5652 13492 -5646
rect 13434 -5686 13446 -5652
rect 13434 -5692 13492 -5686
rect 13434 -5852 13492 -5846
rect 13434 -5886 13446 -5852
rect 13434 -5892 13492 -5886
rect 15100 -5935 15170 -5584
rect 15282 -5652 15340 -5646
rect 15282 -5686 15294 -5652
rect 15282 -5692 15340 -5686
rect 15282 -5852 15340 -5846
rect 15282 -5886 15294 -5852
rect 15282 -5892 15340 -5886
rect 16948 -5935 17018 -5584
rect 17130 -5652 17188 -5646
rect 17130 -5686 17142 -5652
rect 17130 -5692 17188 -5686
rect 17130 -5852 17188 -5846
rect 17130 -5886 17142 -5852
rect 17130 -5892 17188 -5886
rect 18796 -5935 18866 -5584
rect 18978 -5652 19036 -5646
rect 18978 -5686 18990 -5652
rect 18978 -5692 19036 -5686
rect 18978 -5852 19036 -5846
rect 18978 -5886 18990 -5852
rect 18978 -5892 19036 -5886
rect 20644 -5935 20714 -5584
rect 20826 -5652 20884 -5646
rect 20826 -5686 20838 -5652
rect 20826 -5692 20884 -5686
rect 20826 -5852 20884 -5846
rect 20826 -5886 20838 -5852
rect 20826 -5892 20884 -5886
rect 22492 -5935 22562 -5584
rect 22674 -5652 22732 -5646
rect 22674 -5686 22686 -5652
rect 22674 -5692 22732 -5686
rect 22674 -5852 22732 -5846
rect 22674 -5886 22686 -5852
rect 22674 -5892 22732 -5886
rect 24340 -5935 24410 -5584
rect 24522 -5652 24580 -5646
rect 24522 -5686 24534 -5652
rect 24522 -5692 24580 -5686
rect 24522 -5852 24580 -5846
rect 24522 -5886 24534 -5852
rect 24522 -5892 24580 -5886
rect 26188 -5935 26258 -5584
rect 26370 -5652 26428 -5646
rect 26370 -5686 26382 -5652
rect 26370 -5692 26428 -5686
rect 26370 -5852 26428 -5846
rect 26370 -5886 26382 -5852
rect 26370 -5892 26428 -5886
rect 28036 -5935 28106 -5584
rect 28218 -5652 28276 -5646
rect 28218 -5686 28230 -5652
rect 28218 -5692 28276 -5686
rect 28218 -5852 28276 -5846
rect 28218 -5886 28230 -5852
rect 28218 -5892 28276 -5886
rect 29884 -5935 29954 -5584
rect 30066 -5652 30124 -5646
rect 30066 -5686 30078 -5652
rect 30066 -5692 30124 -5686
rect 30066 -5852 30124 -5846
rect 30066 -5886 30078 -5852
rect 30066 -5892 30124 -5886
rect 31732 -5935 31802 -5584
rect 31914 -5652 31972 -5646
rect 31914 -5686 31926 -5652
rect 31914 -5692 31972 -5686
rect 31914 -5852 31972 -5846
rect 31914 -5886 31926 -5852
rect 31914 -5892 31972 -5886
rect 33580 -5935 33650 -5584
rect 33762 -5652 33820 -5646
rect 33762 -5686 33774 -5652
rect 33762 -5692 33820 -5686
rect 33762 -5852 33820 -5846
rect 33762 -5886 33774 -5852
rect 33762 -5892 33820 -5886
rect 35428 -5935 35498 -5584
rect 35610 -5652 35668 -5646
rect 35610 -5686 35622 -5652
rect 35610 -5692 35668 -5686
rect 35610 -5852 35668 -5846
rect 35610 -5886 35622 -5852
rect 35610 -5892 35668 -5886
rect 37276 -5935 37346 -5584
rect 37458 -5652 37516 -5646
rect 37458 -5686 37470 -5652
rect 37458 -5692 37516 -5686
rect 37458 -5852 37516 -5846
rect 37458 -5886 37470 -5852
rect 37458 -5892 37516 -5886
rect 39124 -5935 39194 -5584
rect 39306 -5652 39364 -5646
rect 39306 -5686 39318 -5652
rect 39306 -5692 39364 -5686
rect 39306 -5852 39364 -5846
rect 39306 -5886 39318 -5852
rect 39306 -5892 39364 -5886
rect 40972 -5935 41042 -5584
rect 41154 -5652 41212 -5646
rect 41154 -5686 41166 -5652
rect 41154 -5692 41212 -5686
rect 41154 -5852 41212 -5846
rect 41154 -5886 41166 -5852
rect 41154 -5892 41212 -5886
rect 42820 -5935 42890 -5584
rect 43002 -5652 43060 -5646
rect 43002 -5686 43014 -5652
rect 43002 -5692 43060 -5686
rect 43002 -5852 43060 -5846
rect 43002 -5886 43014 -5852
rect 43002 -5892 43060 -5886
rect 44668 -5935 44738 -5584
rect 44850 -5652 44908 -5646
rect 44850 -5686 44862 -5652
rect 44850 -5692 44908 -5686
rect 44850 -5852 44908 -5846
rect 44850 -5886 44862 -5852
rect 44850 -5892 44908 -5886
rect 46516 -5935 46586 -5584
rect 46698 -5652 46756 -5646
rect 46698 -5686 46710 -5652
rect 46698 -5692 46756 -5686
rect 46698 -5852 46756 -5846
rect 46698 -5886 46710 -5852
rect 46698 -5892 46756 -5886
rect 48364 -5935 48434 -5584
rect 48546 -5652 48604 -5646
rect 48546 -5686 48558 -5652
rect 48546 -5692 48604 -5686
rect 48546 -5852 48604 -5846
rect 48546 -5886 48558 -5852
rect 48546 -5892 48604 -5886
rect 50212 -5935 50282 -5584
rect 50394 -5652 50452 -5646
rect 50394 -5686 50406 -5652
rect 50394 -5692 50452 -5686
rect 50394 -5852 50452 -5846
rect 50394 -5886 50406 -5852
rect 50394 -5892 50452 -5886
rect 52060 -5935 52130 -5584
rect 52242 -5652 52300 -5646
rect 52242 -5686 52254 -5652
rect 52242 -5692 52300 -5686
rect 52242 -5852 52300 -5846
rect 52242 -5886 52254 -5852
rect 52242 -5892 52300 -5886
rect 53908 -5935 53978 -5584
rect 54090 -5652 54148 -5646
rect 54090 -5686 54102 -5652
rect 54090 -5692 54148 -5686
rect 54090 -5852 54148 -5846
rect 54090 -5886 54102 -5852
rect 54090 -5892 54148 -5886
rect 55756 -5935 55826 -5584
rect 55938 -5652 55996 -5646
rect 55938 -5686 55950 -5652
rect 55938 -5692 55996 -5686
rect 55938 -5852 55996 -5846
rect 55938 -5886 55950 -5852
rect 55938 -5892 55996 -5886
rect 57604 -5935 57674 -5584
rect 57786 -5652 57844 -5646
rect 57786 -5686 57798 -5652
rect 57786 -5692 57844 -5686
rect 57786 -5852 57844 -5846
rect 57786 -5886 57798 -5852
rect 57786 -5892 57844 -5886
rect 59452 -5935 59522 -5584
rect 59634 -5652 59692 -5646
rect 59634 -5686 59646 -5652
rect 59634 -5692 59692 -5686
rect 59634 -5852 59692 -5846
rect 59634 -5886 59646 -5852
rect 59634 -5892 59692 -5886
rect 61300 -5935 61370 -5584
rect 61482 -5652 61540 -5646
rect 61482 -5686 61494 -5652
rect 61482 -5692 61540 -5686
rect 61482 -5852 61540 -5846
rect 61482 -5886 61494 -5852
rect 61482 -5892 61540 -5886
rect 63148 -5935 63218 -5584
rect 63330 -5652 63388 -5646
rect 63330 -5686 63342 -5652
rect 63330 -5692 63388 -5686
rect 63330 -5852 63388 -5846
rect 63330 -5886 63342 -5852
rect 63330 -5892 63388 -5886
rect 64996 -5935 65066 -5584
rect 65178 -5652 65236 -5646
rect 65178 -5686 65190 -5652
rect 65178 -5692 65236 -5686
rect 65178 -5852 65236 -5846
rect 65178 -5886 65190 -5852
rect 65178 -5892 65236 -5886
rect 66844 -5935 66914 -5584
rect 67026 -5652 67084 -5646
rect 67026 -5686 67038 -5652
rect 67026 -5692 67084 -5686
rect 67026 -5852 67084 -5846
rect 67026 -5886 67038 -5852
rect 67026 -5892 67084 -5886
rect 68692 -5935 68762 -5584
rect 68874 -5652 68932 -5646
rect 68874 -5686 68886 -5652
rect 68874 -5692 68932 -5686
rect 68874 -5852 68932 -5846
rect 68874 -5886 68886 -5852
rect 68874 -5892 68932 -5886
rect 70540 -5935 70610 -5584
rect 70722 -5652 70780 -5646
rect 70722 -5686 70734 -5652
rect 70722 -5692 70780 -5686
rect 70722 -5852 70780 -5846
rect 70722 -5886 70734 -5852
rect 70722 -5892 70780 -5886
rect 72388 -5935 72458 -5584
rect 72570 -5652 72628 -5646
rect 72570 -5686 72582 -5652
rect 72570 -5692 72628 -5686
rect 72570 -5852 72628 -5846
rect 72570 -5886 72582 -5852
rect 72570 -5892 72628 -5886
rect 74236 -5935 74306 -5584
rect 74418 -5652 74476 -5646
rect 74418 -5686 74430 -5652
rect 74418 -5692 74476 -5686
rect 74418 -5852 74476 -5846
rect 74418 -5886 74430 -5852
rect 74418 -5892 74476 -5886
rect 76084 -5935 76154 -5584
rect 76266 -5652 76324 -5646
rect 76266 -5686 76278 -5652
rect 76266 -5692 76324 -5686
rect 76266 -5852 76324 -5846
rect 76266 -5886 76278 -5852
rect 76266 -5892 76324 -5886
rect 77932 -5935 78002 -5584
rect 78114 -5652 78172 -5646
rect 78114 -5686 78126 -5652
rect 78114 -5692 78172 -5686
rect 78114 -5852 78172 -5846
rect 78114 -5886 78126 -5852
rect 78114 -5892 78172 -5886
rect 79780 -5935 79850 -5584
rect 79962 -5652 80020 -5646
rect 79962 -5686 79974 -5652
rect 79962 -5692 80020 -5686
rect 79962 -5852 80020 -5846
rect 79962 -5886 79974 -5852
rect 79962 -5892 80020 -5886
rect 81628 -5935 81698 -5584
rect 81810 -5652 81868 -5646
rect 81810 -5686 81822 -5652
rect 81810 -5692 81868 -5686
rect 81810 -5852 81868 -5846
rect 81810 -5886 81822 -5852
rect 81810 -5892 81868 -5886
rect 83476 -5935 83546 -5584
rect 83658 -5652 83716 -5646
rect 83658 -5686 83670 -5652
rect 83658 -5692 83716 -5686
rect 83658 -5852 83716 -5846
rect 83658 -5886 83670 -5852
rect 83658 -5892 83716 -5886
rect 85324 -5935 85394 -5584
rect 85506 -5652 85564 -5646
rect 85506 -5686 85518 -5652
rect 85506 -5692 85564 -5686
rect 85506 -5852 85564 -5846
rect 85506 -5886 85518 -5852
rect 85506 -5892 85564 -5886
rect 87172 -5935 87242 -5584
rect 87354 -5652 87412 -5646
rect 87354 -5686 87366 -5652
rect 87354 -5692 87412 -5686
rect 87354 -5852 87412 -5846
rect 87354 -5886 87366 -5852
rect 87354 -5892 87412 -5886
rect 89020 -5935 89090 -5584
rect 89202 -5652 89260 -5646
rect 89202 -5686 89214 -5652
rect 89202 -5692 89260 -5686
rect 89202 -5852 89260 -5846
rect 89202 -5886 89214 -5852
rect 89202 -5892 89260 -5886
rect 90868 -5935 90938 -5584
rect 91050 -5652 91108 -5646
rect 91050 -5686 91062 -5652
rect 91050 -5692 91108 -5686
rect 91050 -5852 91108 -5846
rect 91050 -5886 91062 -5852
rect 91050 -5892 91108 -5886
rect 92716 -5935 92786 -5584
rect 92898 -5652 92956 -5646
rect 92898 -5686 92910 -5652
rect 92898 -5692 92956 -5686
rect 92898 -5852 92956 -5846
rect 92898 -5886 92910 -5852
rect 92898 -5892 92956 -5886
rect 94564 -5935 94634 -5584
rect 94746 -5652 94804 -5646
rect 94746 -5686 94758 -5652
rect 94746 -5692 94804 -5686
rect 94746 -5852 94804 -5846
rect 94746 -5886 94758 -5852
rect 94746 -5892 94804 -5886
rect 96412 -5935 96482 -5584
rect 96594 -5652 96652 -5646
rect 96594 -5686 96606 -5652
rect 96594 -5692 96652 -5686
rect 96594 -5852 96652 -5846
rect 96594 -5886 96606 -5852
rect 96594 -5892 96652 -5886
rect 98260 -5935 98330 -5584
rect 98442 -5652 98500 -5646
rect 98442 -5686 98454 -5652
rect 98442 -5692 98500 -5686
rect 98442 -5852 98500 -5846
rect 98442 -5886 98454 -5852
rect 98442 -5892 98500 -5886
rect 100108 -5935 100178 -5584
rect 100290 -5652 100348 -5646
rect 100290 -5686 100302 -5652
rect 100290 -5692 100348 -5686
rect 100290 -5852 100348 -5846
rect 100290 -5886 100302 -5852
rect 100290 -5892 100348 -5886
rect 101956 -5935 102026 -5584
rect 102138 -5652 102196 -5646
rect 102138 -5686 102150 -5652
rect 102138 -5692 102196 -5686
rect 102138 -5852 102196 -5846
rect 102138 -5886 102150 -5852
rect 102138 -5892 102196 -5886
rect 103804 -5935 103874 -5584
rect 103986 -5652 104044 -5646
rect 103986 -5686 103998 -5652
rect 103986 -5692 104044 -5686
rect 103986 -5852 104044 -5846
rect 103986 -5886 103998 -5852
rect 103986 -5892 104044 -5886
rect 105652 -5935 105722 -5584
rect 105834 -5652 105892 -5646
rect 105834 -5686 105846 -5652
rect 105834 -5692 105892 -5686
rect 105834 -5852 105892 -5846
rect 105834 -5886 105846 -5852
rect 105834 -5892 105892 -5886
rect 107500 -5935 107570 -5584
rect 107682 -5652 107740 -5646
rect 107682 -5686 107694 -5652
rect 107682 -5692 107740 -5686
rect 107682 -5852 107740 -5846
rect 107682 -5886 107694 -5852
rect 107682 -5892 107740 -5886
rect 109348 -5935 109418 -5584
rect 109530 -5652 109588 -5646
rect 109530 -5686 109542 -5652
rect 109530 -5692 109588 -5686
rect 109530 -5852 109588 -5846
rect 109530 -5886 109542 -5852
rect 109530 -5892 109588 -5886
rect 111196 -5935 111266 -5584
rect 111378 -5652 111436 -5646
rect 111378 -5686 111390 -5652
rect 111378 -5692 111436 -5686
rect 111378 -5852 111436 -5846
rect 111378 -5886 111390 -5852
rect 111378 -5892 111436 -5886
rect 113044 -5935 113114 -5584
rect 113226 -5652 113284 -5646
rect 113226 -5686 113238 -5652
rect 113226 -5692 113284 -5686
rect 113226 -5852 113284 -5846
rect 113226 -5886 113238 -5852
rect 113226 -5892 113284 -5886
rect 114892 -5935 114962 -5584
rect 115074 -5652 115132 -5646
rect 115074 -5686 115086 -5652
rect 115074 -5692 115132 -5686
rect 115074 -5852 115132 -5846
rect 115074 -5886 115086 -5852
rect 115074 -5892 115132 -5886
rect 116740 -5935 116810 -5584
rect 116922 -5652 116980 -5646
rect 116922 -5686 116934 -5652
rect 116922 -5692 116980 -5686
rect 116922 -5852 116980 -5846
rect 116922 -5886 116934 -5852
rect 116922 -5892 116980 -5886
rect 118588 -5935 118658 -5584
rect 118770 -5652 118828 -5646
rect 118770 -5686 118782 -5652
rect 118770 -5692 118828 -5686
rect 118770 -5852 118828 -5846
rect 118770 -5886 118782 -5852
rect 118770 -5892 118828 -5886
rect 120436 -5935 120506 -5584
rect 120618 -5652 120676 -5646
rect 120618 -5686 120630 -5652
rect 120618 -5692 120676 -5686
rect 120618 -5852 120676 -5846
rect 120618 -5886 120630 -5852
rect 120618 -5892 120676 -5886
rect 122284 -5935 122354 -5584
rect 122466 -5652 122524 -5646
rect 122466 -5686 122478 -5652
rect 122466 -5692 122524 -5686
rect 122466 -5852 122524 -5846
rect 122466 -5886 122478 -5852
rect 122466 -5892 122524 -5886
rect 124132 -5935 124202 -5584
rect 124314 -5652 124372 -5646
rect 124314 -5686 124326 -5652
rect 124314 -5692 124372 -5686
rect 124314 -5852 124372 -5846
rect 124314 -5886 124326 -5852
rect 124314 -5892 124372 -5886
rect 125980 -5935 126050 -5584
rect 126162 -5652 126220 -5646
rect 126162 -5686 126174 -5652
rect 126162 -5692 126220 -5686
rect 126162 -5852 126220 -5846
rect 126162 -5886 126174 -5852
rect 126162 -5892 126220 -5886
rect 127828 -5935 127898 -5584
rect 128010 -5652 128068 -5646
rect 128010 -5686 128022 -5652
rect 128010 -5692 128068 -5686
rect 128010 -5852 128068 -5846
rect 128010 -5886 128022 -5852
rect 128010 -5892 128068 -5886
rect 129676 -5935 129746 -5584
rect 129858 -5652 129916 -5646
rect 129858 -5686 129870 -5652
rect 129858 -5692 129916 -5686
rect 129858 -5852 129916 -5846
rect 129858 -5886 129870 -5852
rect 129858 -5892 129916 -5886
rect 131524 -5935 131594 -5584
rect 131706 -5652 131764 -5646
rect 131706 -5686 131718 -5652
rect 131706 -5692 131764 -5686
rect 131706 -5852 131764 -5846
rect 131706 -5886 131718 -5852
rect 131706 -5892 131764 -5886
rect 133372 -5935 133442 -5584
rect 133554 -5652 133612 -5646
rect 133554 -5686 133566 -5652
rect 133554 -5692 133612 -5686
rect 133554 -5852 133612 -5846
rect 133554 -5886 133566 -5852
rect 133554 -5892 133612 -5886
rect 135220 -5935 135290 -5584
rect 135402 -5652 135460 -5646
rect 135402 -5686 135414 -5652
rect 135402 -5692 135460 -5686
rect 135402 -5852 135460 -5846
rect 135402 -5886 135414 -5852
rect 135402 -5892 135460 -5886
rect 137068 -5935 137138 -5584
rect 137250 -5652 137308 -5646
rect 137250 -5686 137262 -5652
rect 137250 -5692 137308 -5686
rect 137250 -5852 137308 -5846
rect 137250 -5886 137262 -5852
rect 137250 -5892 137308 -5886
rect 138916 -5935 138986 -5584
rect 139098 -5652 139156 -5646
rect 139098 -5686 139110 -5652
rect 139098 -5692 139156 -5686
rect 139098 -5852 139156 -5846
rect 139098 -5886 139110 -5852
rect 139098 -5892 139156 -5886
rect 140764 -5935 140834 -5584
rect 140946 -5652 141004 -5646
rect 140946 -5686 140958 -5652
rect 140946 -5692 141004 -5686
rect 140946 -5852 141004 -5846
rect 140946 -5886 140958 -5852
rect 140946 -5892 141004 -5886
rect 142612 -5935 142682 -5584
rect 142794 -5652 142852 -5646
rect 142794 -5686 142806 -5652
rect 142794 -5692 142852 -5686
rect 142794 -5852 142852 -5846
rect 142794 -5886 142806 -5852
rect 142794 -5892 142852 -5886
rect 144460 -5935 144530 -5584
rect 144642 -5652 144700 -5646
rect 144642 -5686 144654 -5652
rect 144642 -5692 144700 -5686
rect 144642 -5852 144700 -5846
rect 144642 -5886 144654 -5852
rect 144642 -5892 144700 -5886
rect 146308 -5935 146378 -5584
rect 146490 -5652 146548 -5646
rect 146490 -5686 146502 -5652
rect 146490 -5692 146548 -5686
rect 146490 -5852 146548 -5846
rect 146490 -5886 146502 -5852
rect 146490 -5892 146548 -5886
rect 148156 -5935 148226 -5584
rect 148338 -5652 148396 -5646
rect 148338 -5686 148350 -5652
rect 148338 -5692 148396 -5686
rect 148338 -5852 148396 -5846
rect 148338 -5886 148350 -5852
rect 148338 -5892 148396 -5886
rect 150004 -5935 150074 -5584
rect 150186 -5652 150244 -5646
rect 150186 -5686 150198 -5652
rect 150186 -5692 150244 -5686
rect 150186 -5852 150244 -5846
rect 150186 -5886 150198 -5852
rect 150186 -5892 150244 -5886
rect 151852 -5935 151922 -5584
rect 152034 -5652 152092 -5646
rect 152034 -5686 152046 -5652
rect 152034 -5692 152092 -5686
rect 152034 -5852 152092 -5846
rect 152034 -5886 152046 -5852
rect 152034 -5892 152092 -5886
rect 153700 -5935 153770 -5584
rect 153882 -5652 153940 -5646
rect 153882 -5686 153894 -5652
rect 153882 -5692 153940 -5686
rect 153882 -5852 153940 -5846
rect 153882 -5886 153894 -5852
rect 153882 -5892 153940 -5886
rect 155548 -5935 155618 -5584
rect 155730 -5652 155788 -5646
rect 155730 -5686 155742 -5652
rect 155730 -5692 155788 -5686
rect 155730 -5852 155788 -5846
rect 155730 -5886 155742 -5852
rect 155730 -5892 155788 -5886
rect 157396 -5935 157466 -5584
rect 157578 -5652 157636 -5646
rect 157578 -5686 157590 -5652
rect 157578 -5692 157636 -5686
rect 157578 -5852 157636 -5846
rect 157578 -5886 157590 -5852
rect 157578 -5892 157636 -5886
rect 159244 -5935 159314 -5584
rect 159426 -5652 159484 -5646
rect 159426 -5686 159438 -5652
rect 159426 -5692 159484 -5686
rect 159426 -5852 159484 -5846
rect 159426 -5886 159438 -5852
rect 159426 -5892 159484 -5886
rect 161092 -5935 161162 -5584
rect 161274 -5652 161332 -5646
rect 161274 -5686 161286 -5652
rect 161274 -5692 161332 -5686
rect 161274 -5852 161332 -5846
rect 161274 -5886 161286 -5852
rect 161274 -5892 161332 -5886
rect 162940 -5935 163010 -5584
rect 163122 -5652 163180 -5646
rect 163122 -5686 163134 -5652
rect 163122 -5692 163180 -5686
rect 163122 -5852 163180 -5846
rect 163122 -5886 163134 -5852
rect 163122 -5892 163180 -5886
rect 164788 -5935 164858 -5584
rect 164970 -5652 165028 -5646
rect 164970 -5686 164982 -5652
rect 164970 -5692 165028 -5686
rect 164970 -5852 165028 -5846
rect 164970 -5886 164982 -5852
rect 164970 -5892 165028 -5886
rect 166636 -5935 166706 -5584
rect 166818 -5652 166876 -5646
rect 166818 -5686 166830 -5652
rect 166818 -5692 166876 -5686
rect 166818 -5852 166876 -5846
rect 166818 -5886 166830 -5852
rect 166818 -5892 166876 -5886
rect 168484 -5935 168554 -5584
rect 168666 -5652 168724 -5646
rect 168666 -5686 168678 -5652
rect 168666 -5692 168724 -5686
rect 168666 -5852 168724 -5846
rect 168666 -5886 168678 -5852
rect 168666 -5892 168724 -5886
rect 170332 -5935 170402 -5584
rect 170514 -5652 170572 -5646
rect 170514 -5686 170526 -5652
rect 170514 -5692 170572 -5686
rect 170514 -5852 170572 -5846
rect 170514 -5886 170526 -5852
rect 170514 -5892 170572 -5886
rect 172180 -5935 172250 -5584
rect 172362 -5652 172420 -5646
rect 172362 -5686 172374 -5652
rect 172362 -5692 172420 -5686
rect 172362 -5852 172420 -5846
rect 172362 -5886 172374 -5852
rect 172362 -5892 172420 -5886
rect 174028 -5935 174098 -5584
rect 174210 -5652 174268 -5646
rect 174210 -5686 174222 -5652
rect 174210 -5692 174268 -5686
rect 174210 -5852 174268 -5846
rect 174210 -5886 174222 -5852
rect 174210 -5892 174268 -5886
rect 175876 -5935 175946 -5584
rect 176058 -5652 176116 -5646
rect 176058 -5686 176070 -5652
rect 176058 -5692 176116 -5686
rect 176058 -5852 176116 -5846
rect 176058 -5886 176070 -5852
rect 176058 -5892 176116 -5886
rect 177724 -5935 177794 -5584
rect 179332 -5615 179344 -5581
rect 179519 -5584 179590 -5550
rect 179332 -5621 179390 -5615
rect 177906 -5652 177964 -5646
rect 177906 -5686 177918 -5652
rect 177906 -5692 177964 -5686
rect 177906 -5852 177964 -5846
rect 177906 -5886 177918 -5852
rect 177906 -5892 177964 -5886
rect 179519 -5935 179589 -5584
rect 179701 -5652 179759 -5646
rect 179701 -5686 179713 -5652
rect 179701 -5692 179759 -5686
rect 179701 -5852 179759 -5846
rect 179701 -5886 179713 -5852
rect 179701 -5892 179759 -5886
rect 179888 -5901 179958 -5514
rect 180240 -5514 180274 -5513
rect 180662 -5513 180697 -5496
rect 180977 -5513 181012 -5496
rect 180662 -5514 180696 -5513
rect 180240 -5550 180310 -5514
rect 180070 -5581 180128 -5575
rect 180070 -5615 180082 -5581
rect 180257 -5584 180328 -5550
rect 180070 -5621 180128 -5615
rect 179888 -5935 179959 -5901
rect 180257 -5935 180327 -5584
rect 180439 -5652 180497 -5646
rect 180439 -5686 180451 -5652
rect 180439 -5692 180497 -5686
rect 180439 -5852 180497 -5846
rect 180439 -5886 180451 -5852
rect 180439 -5892 180497 -5886
rect 180626 -5901 180696 -5514
rect 180978 -5514 181012 -5513
rect 181400 -5513 181435 -5496
rect 181715 -5513 181750 -5496
rect 181400 -5514 181434 -5513
rect 180978 -5550 181048 -5514
rect 180808 -5581 180866 -5575
rect 180808 -5615 180820 -5581
rect 180995 -5584 181066 -5550
rect 180808 -5621 180866 -5615
rect 180626 -5935 180697 -5901
rect 180995 -5935 181065 -5584
rect 181177 -5652 181235 -5646
rect 181177 -5686 181189 -5652
rect 181177 -5692 181235 -5686
rect 181177 -5852 181235 -5846
rect 181177 -5886 181189 -5852
rect 181177 -5892 181235 -5886
rect 181364 -5901 181434 -5514
rect 181716 -5514 181750 -5513
rect 182138 -5513 182173 -5496
rect 182453 -5513 182488 -5496
rect 182138 -5514 182172 -5513
rect 181716 -5550 181786 -5514
rect 181546 -5581 181604 -5575
rect 181546 -5615 181558 -5581
rect 181733 -5584 181804 -5550
rect 181546 -5621 181604 -5615
rect 181364 -5935 181435 -5901
rect 181733 -5935 181803 -5584
rect 181915 -5652 181973 -5646
rect 181915 -5686 181927 -5652
rect 181915 -5692 181973 -5686
rect 181915 -5852 181973 -5846
rect 181915 -5886 181927 -5852
rect 181915 -5892 181973 -5886
rect 182102 -5901 182172 -5514
rect 182454 -5514 182488 -5513
rect 182876 -5513 182911 -5496
rect 183191 -5513 183226 -5496
rect 182876 -5514 182910 -5513
rect 182454 -5550 182524 -5514
rect 182284 -5581 182342 -5575
rect 182284 -5615 182296 -5581
rect 182471 -5584 182542 -5550
rect 182284 -5621 182342 -5615
rect 182102 -5935 182173 -5901
rect 182471 -5935 182541 -5584
rect 182653 -5652 182711 -5646
rect 182653 -5686 182665 -5652
rect 182653 -5692 182711 -5686
rect 182653 -5852 182711 -5846
rect 182653 -5886 182665 -5852
rect 182653 -5892 182711 -5886
rect 182840 -5901 182910 -5514
rect 183192 -5514 183226 -5513
rect 183614 -5513 183649 -5496
rect 183929 -5513 183964 -5496
rect 183614 -5514 183648 -5513
rect 183192 -5550 183262 -5514
rect 183022 -5581 183080 -5575
rect 183022 -5615 183034 -5581
rect 183209 -5584 183280 -5550
rect 183022 -5621 183080 -5615
rect 182840 -5935 182911 -5901
rect 183209 -5935 183279 -5584
rect 183391 -5652 183449 -5646
rect 183391 -5686 183403 -5652
rect 183391 -5692 183449 -5686
rect 183391 -5852 183449 -5846
rect 183391 -5886 183403 -5852
rect 183391 -5892 183449 -5886
rect 183578 -5901 183648 -5514
rect 183930 -5514 183964 -5513
rect 184352 -5513 184387 -5496
rect 184667 -5513 184702 -5496
rect 184352 -5514 184386 -5513
rect 183930 -5550 184000 -5514
rect 183760 -5581 183818 -5575
rect 183760 -5615 183772 -5581
rect 183947 -5584 184018 -5550
rect 183760 -5621 183818 -5615
rect 183578 -5935 183649 -5901
rect 183947 -5935 184017 -5584
rect 184129 -5652 184187 -5646
rect 184129 -5686 184141 -5652
rect 184129 -5692 184187 -5686
rect 184129 -5852 184187 -5846
rect 184129 -5886 184141 -5852
rect 184129 -5892 184187 -5886
rect 184316 -5901 184386 -5514
rect 184668 -5514 184702 -5513
rect 185090 -5513 185125 -5496
rect 185405 -5513 185440 -5496
rect 185090 -5514 185124 -5513
rect 184668 -5550 184738 -5514
rect 184498 -5581 184556 -5575
rect 184498 -5615 184510 -5581
rect 184685 -5584 184756 -5550
rect 184498 -5621 184556 -5615
rect 184316 -5935 184387 -5901
rect 184685 -5935 184755 -5584
rect 184867 -5652 184925 -5646
rect 184867 -5686 184879 -5652
rect 184867 -5692 184925 -5686
rect 184867 -5852 184925 -5846
rect 184867 -5886 184879 -5852
rect 184867 -5892 184925 -5886
rect 185054 -5901 185124 -5514
rect 185406 -5514 185440 -5513
rect 185828 -5513 185863 -5496
rect 186143 -5513 186178 -5496
rect 185828 -5514 185862 -5513
rect 185406 -5550 185476 -5514
rect 185236 -5581 185294 -5575
rect 185236 -5615 185248 -5581
rect 185423 -5584 185494 -5550
rect 185236 -5621 185294 -5615
rect 185054 -5935 185125 -5901
rect 185423 -5935 185493 -5584
rect 185605 -5652 185663 -5646
rect 185605 -5686 185617 -5652
rect 185605 -5692 185663 -5686
rect 185605 -5852 185663 -5846
rect 185605 -5886 185617 -5852
rect 185605 -5892 185663 -5886
rect 185792 -5901 185862 -5514
rect 186144 -5514 186178 -5513
rect 186566 -5513 186601 -5496
rect 186881 -5513 186916 -5496
rect 186566 -5514 186600 -5513
rect 186144 -5550 186214 -5514
rect 185974 -5581 186032 -5575
rect 185974 -5615 185986 -5581
rect 186161 -5584 186232 -5550
rect 185974 -5621 186032 -5615
rect 185792 -5935 185863 -5901
rect 186161 -5935 186231 -5584
rect 186343 -5652 186401 -5646
rect 186343 -5686 186355 -5652
rect 186343 -5692 186401 -5686
rect 186343 -5852 186401 -5846
rect 186343 -5886 186355 -5852
rect 186343 -5892 186401 -5886
rect 186530 -5901 186600 -5514
rect 186882 -5514 186916 -5513
rect 187304 -5513 187339 -5496
rect 187619 -5513 187654 -5496
rect 187304 -5514 187338 -5513
rect 186882 -5550 186952 -5514
rect 186712 -5581 186770 -5575
rect 186712 -5615 186724 -5581
rect 186899 -5584 186970 -5550
rect 186712 -5621 186770 -5615
rect 186530 -5935 186601 -5901
rect 186899 -5935 186969 -5584
rect 187081 -5652 187139 -5646
rect 187081 -5686 187093 -5652
rect 187081 -5692 187139 -5686
rect 187081 -5852 187139 -5846
rect 187081 -5886 187093 -5852
rect 187081 -5892 187139 -5886
rect 187268 -5901 187338 -5514
rect 187620 -5514 187654 -5513
rect 188042 -5513 188077 -5496
rect 188357 -5513 188392 -5496
rect 188042 -5514 188076 -5513
rect 187620 -5550 187690 -5514
rect 187450 -5581 187508 -5575
rect 187450 -5615 187462 -5581
rect 187637 -5584 187708 -5550
rect 187450 -5621 187508 -5615
rect 187268 -5935 187339 -5901
rect 187637 -5935 187707 -5584
rect 187819 -5652 187877 -5646
rect 187819 -5686 187831 -5652
rect 187819 -5692 187877 -5686
rect 187819 -5852 187877 -5846
rect 187819 -5886 187831 -5852
rect 187819 -5892 187877 -5886
rect 188006 -5901 188076 -5514
rect 188358 -5514 188392 -5513
rect 188780 -5513 188815 -5496
rect 189095 -5513 189130 -5496
rect 188780 -5514 188814 -5513
rect 188358 -5550 188428 -5514
rect 188188 -5581 188246 -5575
rect 188188 -5615 188200 -5581
rect 188375 -5584 188446 -5550
rect 188188 -5621 188246 -5615
rect 188006 -5935 188077 -5901
rect 188375 -5935 188445 -5584
rect 188557 -5652 188615 -5646
rect 188557 -5686 188569 -5652
rect 188557 -5692 188615 -5686
rect 188557 -5852 188615 -5846
rect 188557 -5886 188569 -5852
rect 188557 -5892 188615 -5886
rect 188744 -5901 188814 -5514
rect 189096 -5514 189130 -5513
rect 189518 -5513 189553 -5496
rect 189833 -5513 189868 -5496
rect 189518 -5514 189552 -5513
rect 189096 -5550 189166 -5514
rect 188926 -5581 188984 -5575
rect 188926 -5615 188938 -5581
rect 189113 -5584 189184 -5550
rect 188926 -5621 188984 -5615
rect 188744 -5935 188815 -5901
rect 189113 -5935 189183 -5584
rect 189295 -5652 189353 -5646
rect 189295 -5686 189307 -5652
rect 189295 -5692 189353 -5686
rect 189295 -5852 189353 -5846
rect 189295 -5886 189307 -5852
rect 189295 -5892 189353 -5886
rect 189482 -5901 189552 -5514
rect 189834 -5514 189868 -5513
rect 190256 -5513 190291 -5496
rect 190571 -5513 190606 -5496
rect 190256 -5514 190290 -5513
rect 189834 -5550 189904 -5514
rect 189664 -5581 189722 -5575
rect 189664 -5615 189676 -5581
rect 189851 -5584 189922 -5550
rect 189664 -5621 189722 -5615
rect 189482 -5935 189553 -5901
rect 189851 -5935 189921 -5584
rect 190033 -5652 190091 -5646
rect 190033 -5686 190045 -5652
rect 190033 -5692 190091 -5686
rect 190033 -5852 190091 -5846
rect 190033 -5886 190045 -5852
rect 190033 -5892 190091 -5886
rect 190220 -5901 190290 -5514
rect 190572 -5514 190606 -5513
rect 190994 -5513 191029 -5496
rect 191309 -5513 191344 -5496
rect 190994 -5514 191028 -5513
rect 190572 -5550 190642 -5514
rect 190402 -5581 190460 -5575
rect 190402 -5615 190414 -5581
rect 190589 -5584 190660 -5550
rect 190402 -5621 190460 -5615
rect 190220 -5935 190291 -5901
rect 190589 -5935 190659 -5584
rect 190771 -5652 190829 -5646
rect 190771 -5686 190783 -5652
rect 190771 -5692 190829 -5686
rect 190771 -5852 190829 -5846
rect 190771 -5886 190783 -5852
rect 190771 -5892 190829 -5886
rect 190958 -5901 191028 -5514
rect 191310 -5514 191344 -5513
rect 191732 -5513 191767 -5496
rect 192047 -5513 192082 -5496
rect 191732 -5514 191766 -5513
rect 191310 -5550 191380 -5514
rect 191140 -5581 191198 -5575
rect 191140 -5615 191152 -5581
rect 191327 -5584 191398 -5550
rect 191140 -5621 191198 -5615
rect 190958 -5935 191029 -5901
rect 191327 -5935 191397 -5584
rect 191509 -5652 191567 -5646
rect 191509 -5686 191521 -5652
rect 191509 -5692 191567 -5686
rect 191509 -5852 191567 -5846
rect 191509 -5886 191521 -5852
rect 191509 -5892 191567 -5886
rect 191696 -5901 191766 -5514
rect 192048 -5514 192082 -5513
rect 192470 -5513 192505 -5496
rect 192785 -5513 192820 -5496
rect 192470 -5514 192504 -5513
rect 192048 -5550 192118 -5514
rect 191878 -5581 191936 -5575
rect 191878 -5615 191890 -5581
rect 192065 -5584 192136 -5550
rect 191878 -5621 191936 -5615
rect 191696 -5935 191767 -5901
rect 192065 -5935 192135 -5584
rect 192247 -5652 192305 -5646
rect 192247 -5686 192259 -5652
rect 192247 -5692 192305 -5686
rect 192247 -5852 192305 -5846
rect 192247 -5886 192259 -5852
rect 192247 -5892 192305 -5886
rect 192434 -5901 192504 -5514
rect 192786 -5514 192820 -5513
rect 193208 -5513 193243 -5496
rect 193523 -5513 193558 -5496
rect 193208 -5514 193242 -5513
rect 192786 -5550 192856 -5514
rect 192616 -5581 192674 -5575
rect 192616 -5615 192628 -5581
rect 192803 -5584 192874 -5550
rect 192616 -5621 192674 -5615
rect 192434 -5935 192505 -5901
rect 192803 -5935 192873 -5584
rect 192985 -5652 193043 -5646
rect 192985 -5686 192997 -5652
rect 192985 -5692 193043 -5686
rect 192985 -5852 193043 -5846
rect 192985 -5886 192997 -5852
rect 192985 -5892 193043 -5886
rect 193172 -5901 193242 -5514
rect 193524 -5514 193558 -5513
rect 193946 -5513 193981 -5496
rect 194261 -5513 194296 -5496
rect 193946 -5514 193980 -5513
rect 193524 -5550 193594 -5514
rect 193354 -5581 193412 -5575
rect 193354 -5615 193366 -5581
rect 193541 -5584 193612 -5550
rect 193354 -5621 193412 -5615
rect 193172 -5935 193243 -5901
rect 193541 -5935 193611 -5584
rect 193723 -5652 193781 -5646
rect 193723 -5686 193735 -5652
rect 193723 -5692 193781 -5686
rect 193723 -5852 193781 -5846
rect 193723 -5886 193735 -5852
rect 193723 -5892 193781 -5886
rect 193910 -5901 193980 -5514
rect 194262 -5514 194296 -5513
rect 194684 -5513 194719 -5496
rect 194999 -5513 195034 -5496
rect 194684 -5514 194718 -5513
rect 194262 -5550 194332 -5514
rect 194092 -5581 194150 -5575
rect 194092 -5615 194104 -5581
rect 194279 -5584 194350 -5550
rect 194092 -5621 194150 -5615
rect 193910 -5935 193981 -5901
rect 194279 -5935 194349 -5584
rect 194461 -5652 194519 -5646
rect 194461 -5686 194473 -5652
rect 194461 -5692 194519 -5686
rect 194461 -5852 194519 -5846
rect 194461 -5886 194473 -5852
rect 194461 -5892 194519 -5886
rect 194648 -5901 194718 -5514
rect 195000 -5514 195034 -5513
rect 195422 -5513 195457 -5496
rect 195737 -5513 195772 -5496
rect 195422 -5514 195456 -5513
rect 195000 -5550 195070 -5514
rect 194830 -5581 194888 -5575
rect 194830 -5615 194842 -5581
rect 195017 -5584 195088 -5550
rect 194830 -5621 194888 -5615
rect 194648 -5935 194719 -5901
rect 195017 -5935 195087 -5584
rect 195199 -5652 195257 -5646
rect 195199 -5686 195211 -5652
rect 195199 -5692 195257 -5686
rect 195199 -5852 195257 -5846
rect 195199 -5886 195211 -5852
rect 195199 -5892 195257 -5886
rect 195386 -5901 195456 -5514
rect 195738 -5514 195772 -5513
rect 196160 -5513 196195 -5496
rect 196475 -5513 196510 -5496
rect 196160 -5514 196194 -5513
rect 195738 -5550 195808 -5514
rect 195568 -5581 195626 -5575
rect 195568 -5615 195580 -5581
rect 195755 -5584 195826 -5550
rect 195568 -5621 195626 -5615
rect 195386 -5935 195457 -5901
rect 195755 -5935 195825 -5584
rect 195937 -5652 195995 -5646
rect 195937 -5686 195949 -5652
rect 195937 -5692 195995 -5686
rect 195937 -5852 195995 -5846
rect 195937 -5886 195949 -5852
rect 195937 -5892 195995 -5886
rect 196124 -5901 196194 -5514
rect 196476 -5514 196510 -5513
rect 196898 -5513 196933 -5496
rect 197213 -5513 197248 -5496
rect 196898 -5514 196932 -5513
rect 196476 -5550 196546 -5514
rect 196306 -5581 196364 -5575
rect 196306 -5615 196318 -5581
rect 196493 -5584 196564 -5550
rect 196306 -5621 196364 -5615
rect 196124 -5935 196195 -5901
rect 196493 -5935 196563 -5584
rect 196675 -5652 196733 -5646
rect 196675 -5686 196687 -5652
rect 196675 -5692 196733 -5686
rect 196675 -5852 196733 -5846
rect 196675 -5886 196687 -5852
rect 196675 -5892 196733 -5886
rect 196862 -5901 196932 -5514
rect 197214 -5514 197248 -5513
rect 197636 -5513 197671 -5496
rect 197951 -5513 197986 -5496
rect 197636 -5514 197670 -5513
rect 197214 -5550 197284 -5514
rect 197044 -5581 197102 -5575
rect 197044 -5615 197056 -5581
rect 197231 -5584 197302 -5550
rect 197044 -5621 197102 -5615
rect 196862 -5935 196933 -5901
rect 197231 -5935 197301 -5584
rect 197413 -5652 197471 -5646
rect 197413 -5686 197425 -5652
rect 197413 -5692 197471 -5686
rect 197413 -5852 197471 -5846
rect 197413 -5886 197425 -5852
rect 197413 -5892 197471 -5886
rect 197600 -5901 197670 -5514
rect 197952 -5514 197986 -5513
rect 198374 -5513 198409 -5496
rect 198689 -5513 198724 -5496
rect 198374 -5514 198408 -5513
rect 197952 -5550 198022 -5514
rect 197782 -5581 197840 -5575
rect 197782 -5615 197794 -5581
rect 197969 -5584 198040 -5550
rect 197782 -5621 197840 -5615
rect 197600 -5935 197671 -5901
rect 197969 -5935 198039 -5584
rect 198151 -5652 198209 -5646
rect 198151 -5686 198163 -5652
rect 198151 -5692 198209 -5686
rect 198151 -5852 198209 -5846
rect 198151 -5886 198163 -5852
rect 198151 -5892 198209 -5886
rect 198338 -5901 198408 -5514
rect 198690 -5514 198724 -5513
rect 199112 -5513 199147 -5496
rect 199427 -5513 199462 -5496
rect 199112 -5514 199146 -5513
rect 198690 -5550 198760 -5514
rect 198520 -5581 198578 -5575
rect 198520 -5615 198532 -5581
rect 198707 -5584 198778 -5550
rect 198520 -5621 198578 -5615
rect 198338 -5935 198409 -5901
rect 198707 -5935 198777 -5584
rect 198889 -5652 198947 -5646
rect 198889 -5686 198901 -5652
rect 198889 -5692 198947 -5686
rect 198889 -5852 198947 -5846
rect 198889 -5886 198901 -5852
rect 198889 -5892 198947 -5886
rect 199076 -5901 199146 -5514
rect 199428 -5514 199462 -5513
rect 199850 -5513 199885 -5496
rect 200165 -5513 200200 -5496
rect 199850 -5514 199884 -5513
rect 199428 -5550 199498 -5514
rect 199258 -5581 199316 -5575
rect 199258 -5615 199270 -5581
rect 199445 -5584 199516 -5550
rect 199258 -5621 199316 -5615
rect 199076 -5935 199147 -5901
rect 199445 -5935 199515 -5584
rect 199627 -5652 199685 -5646
rect 199627 -5686 199639 -5652
rect 199627 -5692 199685 -5686
rect 199627 -5852 199685 -5846
rect 199627 -5886 199639 -5852
rect 199627 -5892 199685 -5886
rect 199814 -5901 199884 -5514
rect 200166 -5514 200200 -5513
rect 200588 -5513 200623 -5496
rect 200903 -5513 200938 -5496
rect 200588 -5514 200622 -5513
rect 200166 -5550 200236 -5514
rect 199996 -5581 200054 -5575
rect 199996 -5615 200008 -5581
rect 200183 -5584 200254 -5550
rect 199996 -5621 200054 -5615
rect 199814 -5935 199885 -5901
rect 200183 -5935 200253 -5584
rect 200365 -5652 200423 -5646
rect 200365 -5686 200377 -5652
rect 200365 -5692 200423 -5686
rect 200365 -5852 200423 -5846
rect 200365 -5886 200377 -5852
rect 200365 -5892 200423 -5886
rect 200552 -5901 200622 -5514
rect 200904 -5514 200938 -5513
rect 201326 -5513 201361 -5496
rect 201641 -5513 201676 -5496
rect 201326 -5514 201360 -5513
rect 200904 -5550 200974 -5514
rect 200734 -5581 200792 -5575
rect 200734 -5615 200746 -5581
rect 200921 -5584 200992 -5550
rect 200734 -5621 200792 -5615
rect 200552 -5935 200623 -5901
rect 200921 -5935 200991 -5584
rect 201103 -5652 201161 -5646
rect 201103 -5686 201115 -5652
rect 201103 -5692 201161 -5686
rect 201103 -5852 201161 -5846
rect 201103 -5886 201115 -5852
rect 201103 -5892 201161 -5886
rect 201290 -5901 201360 -5514
rect 201642 -5514 201676 -5513
rect 202064 -5513 202099 -5496
rect 202379 -5513 202414 -5496
rect 202064 -5514 202098 -5513
rect 201642 -5550 201712 -5514
rect 201472 -5581 201530 -5575
rect 201472 -5615 201484 -5581
rect 201659 -5584 201730 -5550
rect 201472 -5621 201530 -5615
rect 201290 -5935 201361 -5901
rect 201659 -5935 201729 -5584
rect 201841 -5652 201899 -5646
rect 201841 -5686 201853 -5652
rect 201841 -5692 201899 -5686
rect 201841 -5852 201899 -5846
rect 201841 -5886 201853 -5852
rect 201841 -5892 201899 -5886
rect 202028 -5901 202098 -5514
rect 202380 -5514 202414 -5513
rect 202802 -5513 202837 -5496
rect 203117 -5513 203152 -5496
rect 202802 -5514 202836 -5513
rect 202380 -5550 202450 -5514
rect 202210 -5581 202268 -5575
rect 202210 -5615 202222 -5581
rect 202397 -5584 202468 -5550
rect 202210 -5621 202268 -5615
rect 202028 -5935 202099 -5901
rect 202397 -5935 202467 -5584
rect 202579 -5652 202637 -5646
rect 202579 -5686 202591 -5652
rect 202579 -5692 202637 -5686
rect 202579 -5852 202637 -5846
rect 202579 -5886 202591 -5852
rect 202579 -5892 202637 -5886
rect 202766 -5901 202836 -5514
rect 203118 -5514 203152 -5513
rect 203540 -5513 203575 -5496
rect 203855 -5513 203890 -5496
rect 203540 -5514 203574 -5513
rect 203118 -5550 203188 -5514
rect 202948 -5581 203006 -5575
rect 202948 -5615 202960 -5581
rect 203135 -5584 203206 -5550
rect 202948 -5621 203006 -5615
rect 202766 -5935 202837 -5901
rect 203135 -5935 203205 -5584
rect 203317 -5652 203375 -5646
rect 203317 -5686 203329 -5652
rect 203317 -5692 203375 -5686
rect 203317 -5852 203375 -5846
rect 203317 -5886 203329 -5852
rect 203317 -5892 203375 -5886
rect 203504 -5901 203574 -5514
rect 203856 -5514 203890 -5513
rect 204278 -5513 204313 -5496
rect 204593 -5513 204628 -5496
rect 204278 -5514 204312 -5513
rect 203856 -5550 203926 -5514
rect 203686 -5581 203744 -5575
rect 203686 -5615 203698 -5581
rect 203873 -5584 203944 -5550
rect 203686 -5621 203744 -5615
rect 203504 -5935 203575 -5901
rect 203873 -5935 203943 -5584
rect 204055 -5652 204113 -5646
rect 204055 -5686 204067 -5652
rect 204055 -5692 204113 -5686
rect 204055 -5852 204113 -5846
rect 204055 -5886 204067 -5852
rect 204055 -5892 204113 -5886
rect 204242 -5901 204312 -5514
rect 204594 -5514 204628 -5513
rect 205016 -5513 205051 -5496
rect 205331 -5513 205366 -5496
rect 205016 -5514 205050 -5513
rect 204594 -5550 204664 -5514
rect 204424 -5581 204482 -5575
rect 204424 -5615 204436 -5581
rect 204611 -5584 204682 -5550
rect 204424 -5621 204482 -5615
rect 204242 -5935 204313 -5901
rect 204611 -5935 204681 -5584
rect 204793 -5652 204851 -5646
rect 204793 -5686 204805 -5652
rect 204793 -5692 204851 -5686
rect 204793 -5852 204851 -5846
rect 204793 -5886 204805 -5852
rect 204793 -5892 204851 -5886
rect 204980 -5901 205050 -5514
rect 205332 -5514 205366 -5513
rect 205754 -5513 205789 -5496
rect 206069 -5513 206104 -5496
rect 205754 -5514 205788 -5513
rect 205332 -5550 205402 -5514
rect 205162 -5581 205220 -5575
rect 205162 -5615 205174 -5581
rect 205349 -5584 205420 -5550
rect 205162 -5621 205220 -5615
rect 204980 -5935 205051 -5901
rect 205349 -5935 205419 -5584
rect 205531 -5652 205589 -5646
rect 205531 -5686 205543 -5652
rect 205531 -5692 205589 -5686
rect 205531 -5852 205589 -5846
rect 205531 -5886 205543 -5852
rect 205531 -5892 205589 -5886
rect 205718 -5901 205788 -5514
rect 206070 -5514 206104 -5513
rect 206492 -5513 206527 -5496
rect 206807 -5513 206842 -5496
rect 206492 -5514 206526 -5513
rect 206070 -5550 206140 -5514
rect 205900 -5581 205958 -5575
rect 205900 -5615 205912 -5581
rect 206087 -5584 206158 -5550
rect 205900 -5621 205958 -5615
rect 205718 -5935 205789 -5901
rect 206087 -5935 206157 -5584
rect 206269 -5652 206327 -5646
rect 206269 -5686 206281 -5652
rect 206269 -5692 206327 -5686
rect 206269 -5852 206327 -5846
rect 206269 -5886 206281 -5852
rect 206269 -5892 206327 -5886
rect 206456 -5901 206526 -5514
rect 206808 -5514 206842 -5513
rect 207230 -5513 207265 -5496
rect 207545 -5513 207580 -5496
rect 207230 -5514 207264 -5513
rect 206808 -5550 206878 -5514
rect 206638 -5581 206696 -5575
rect 206638 -5615 206650 -5581
rect 206825 -5584 206896 -5550
rect 206638 -5621 206696 -5615
rect 206456 -5935 206527 -5901
rect 206825 -5935 206895 -5584
rect 207007 -5652 207065 -5646
rect 207007 -5686 207019 -5652
rect 207007 -5692 207065 -5686
rect 207007 -5852 207065 -5846
rect 207007 -5886 207019 -5852
rect 207007 -5892 207065 -5886
rect 207194 -5901 207264 -5514
rect 207546 -5514 207580 -5513
rect 207968 -5513 208003 -5496
rect 208283 -5513 208318 -5496
rect 207968 -5514 208002 -5513
rect 207546 -5550 207616 -5514
rect 207376 -5581 207434 -5575
rect 207376 -5615 207388 -5581
rect 207563 -5584 207634 -5550
rect 207376 -5621 207434 -5615
rect 207194 -5935 207265 -5901
rect 207563 -5935 207633 -5584
rect 207745 -5652 207803 -5646
rect 207745 -5686 207757 -5652
rect 207745 -5692 207803 -5686
rect 207745 -5852 207803 -5846
rect 207745 -5886 207757 -5852
rect 207745 -5892 207803 -5886
rect 207932 -5901 208002 -5514
rect 208284 -5514 208318 -5513
rect 208706 -5513 208741 -5496
rect 209021 -5513 209056 -5496
rect 208706 -5514 208740 -5513
rect 208284 -5550 208354 -5514
rect 208114 -5581 208172 -5575
rect 208114 -5615 208126 -5581
rect 208301 -5584 208372 -5550
rect 208114 -5621 208172 -5615
rect 207932 -5935 208003 -5901
rect 208301 -5935 208371 -5584
rect 208483 -5652 208541 -5646
rect 208483 -5686 208495 -5652
rect 208483 -5692 208541 -5686
rect 208483 -5852 208541 -5846
rect 208483 -5886 208495 -5852
rect 208483 -5892 208541 -5886
rect 208670 -5901 208740 -5514
rect 209022 -5514 209056 -5513
rect 209444 -5513 209479 -5496
rect 209759 -5513 209794 -5496
rect 209444 -5514 209478 -5513
rect 209022 -5550 209092 -5514
rect 208852 -5581 208910 -5575
rect 208852 -5615 208864 -5581
rect 209039 -5584 209110 -5550
rect 208852 -5621 208910 -5615
rect 208670 -5935 208741 -5901
rect 209039 -5935 209109 -5584
rect 209221 -5652 209279 -5646
rect 209221 -5686 209233 -5652
rect 209221 -5692 209279 -5686
rect 209221 -5852 209279 -5846
rect 209221 -5886 209233 -5852
rect 209221 -5892 209279 -5886
rect 209408 -5901 209478 -5514
rect 209760 -5514 209794 -5513
rect 210182 -5513 210217 -5496
rect 210497 -5513 210532 -5496
rect 210182 -5514 210216 -5513
rect 209760 -5550 209830 -5514
rect 209590 -5581 209648 -5575
rect 209590 -5615 209602 -5581
rect 209777 -5584 209848 -5550
rect 209590 -5621 209648 -5615
rect 209408 -5935 209479 -5901
rect 209777 -5935 209847 -5584
rect 209959 -5652 210017 -5646
rect 209959 -5686 209971 -5652
rect 209959 -5692 210017 -5686
rect 209959 -5852 210017 -5846
rect 209959 -5886 209971 -5852
rect 209959 -5892 210017 -5886
rect 210146 -5901 210216 -5514
rect 210498 -5514 210532 -5513
rect 210920 -5513 210955 -5496
rect 211235 -5513 211270 -5496
rect 210920 -5514 210954 -5513
rect 210498 -5550 210568 -5514
rect 210328 -5581 210386 -5575
rect 210328 -5615 210340 -5581
rect 210515 -5584 210586 -5550
rect 210328 -5621 210386 -5615
rect 210146 -5935 210217 -5901
rect 210515 -5935 210585 -5584
rect 210697 -5652 210755 -5646
rect 210697 -5686 210709 -5652
rect 210697 -5692 210755 -5686
rect 210697 -5852 210755 -5846
rect 210697 -5886 210709 -5852
rect 210697 -5892 210755 -5886
rect 210884 -5901 210954 -5514
rect 211236 -5514 211270 -5513
rect 211658 -5513 211693 -5496
rect 211973 -5513 212008 -5496
rect 211658 -5514 211692 -5513
rect 211236 -5550 211306 -5514
rect 211066 -5581 211124 -5575
rect 211066 -5615 211078 -5581
rect 211253 -5584 211324 -5550
rect 211066 -5621 211124 -5615
rect 210884 -5935 210955 -5901
rect 211253 -5935 211323 -5584
rect 211435 -5652 211493 -5646
rect 211435 -5686 211447 -5652
rect 211435 -5692 211493 -5686
rect 211435 -5852 211493 -5846
rect 211435 -5886 211447 -5852
rect 211435 -5892 211493 -5886
rect 211622 -5901 211692 -5514
rect 211974 -5514 212008 -5513
rect 212396 -5513 212431 -5496
rect 212711 -5513 212746 -5496
rect 212396 -5514 212430 -5513
rect 211974 -5550 212044 -5514
rect 211804 -5581 211862 -5575
rect 211804 -5615 211816 -5581
rect 211991 -5584 212062 -5550
rect 211804 -5621 211862 -5615
rect 211622 -5935 211693 -5901
rect 211991 -5935 212061 -5584
rect 212173 -5652 212231 -5646
rect 212173 -5686 212185 -5652
rect 212173 -5692 212231 -5686
rect 212173 -5852 212231 -5846
rect 212173 -5886 212185 -5852
rect 212173 -5892 212231 -5886
rect 212360 -5901 212430 -5514
rect 212712 -5514 212746 -5513
rect 213134 -5513 213169 -5496
rect 213449 -5513 213484 -5496
rect 213134 -5514 213168 -5513
rect 212712 -5550 212782 -5514
rect 212542 -5581 212600 -5575
rect 212542 -5615 212554 -5581
rect 212729 -5584 212800 -5550
rect 212542 -5621 212600 -5615
rect 212360 -5935 212431 -5901
rect 212729 -5935 212799 -5584
rect 212911 -5652 212969 -5646
rect 212911 -5686 212923 -5652
rect 212911 -5692 212969 -5686
rect 212911 -5852 212969 -5846
rect 212911 -5886 212923 -5852
rect 212911 -5892 212969 -5886
rect 213098 -5901 213168 -5514
rect 213450 -5514 213484 -5513
rect 213872 -5513 213907 -5496
rect 214187 -5513 214222 -5496
rect 213872 -5514 213906 -5513
rect 213450 -5550 213520 -5514
rect 213280 -5581 213338 -5575
rect 213280 -5615 213292 -5581
rect 213467 -5584 213538 -5550
rect 213280 -5621 213338 -5615
rect 213098 -5935 213169 -5901
rect 213467 -5935 213537 -5584
rect 213649 -5652 213707 -5646
rect 213649 -5686 213661 -5652
rect 213649 -5692 213707 -5686
rect 213649 -5852 213707 -5846
rect 213649 -5886 213661 -5852
rect 213649 -5892 213707 -5886
rect 213836 -5901 213906 -5514
rect 214188 -5514 214222 -5513
rect 214610 -5513 214645 -5496
rect 214925 -5513 214960 -5496
rect 214610 -5514 214644 -5513
rect 214188 -5550 214258 -5514
rect 214018 -5581 214076 -5575
rect 214018 -5615 214030 -5581
rect 214205 -5584 214276 -5550
rect 214018 -5621 214076 -5615
rect 213836 -5935 213907 -5901
rect 214205 -5935 214275 -5584
rect 214387 -5652 214445 -5646
rect 214387 -5686 214399 -5652
rect 214387 -5692 214445 -5686
rect 214387 -5852 214445 -5846
rect 214387 -5886 214399 -5852
rect 214387 -5892 214445 -5886
rect 214574 -5901 214644 -5514
rect 214926 -5514 214960 -5513
rect 215348 -5513 215383 -5496
rect 215663 -5513 215698 -5496
rect 215348 -5514 215382 -5513
rect 214926 -5550 214996 -5514
rect 214756 -5581 214814 -5575
rect 214756 -5615 214768 -5581
rect 214943 -5584 215014 -5550
rect 214756 -5621 214814 -5615
rect 214574 -5935 214645 -5901
rect 214943 -5935 215013 -5584
rect 215125 -5652 215183 -5646
rect 215125 -5686 215137 -5652
rect 215125 -5692 215183 -5686
rect 215125 -5852 215183 -5846
rect 215125 -5886 215137 -5852
rect 215125 -5892 215183 -5886
rect 215312 -5901 215382 -5514
rect 215664 -5514 215698 -5513
rect 216086 -5513 216121 -5496
rect 216401 -5513 216436 -5496
rect 216086 -5514 216120 -5513
rect 215664 -5550 215734 -5514
rect 215494 -5581 215552 -5575
rect 215494 -5615 215506 -5581
rect 215681 -5584 215752 -5550
rect 215494 -5621 215552 -5615
rect 215312 -5935 215383 -5901
rect 215681 -5935 215751 -5584
rect 215863 -5652 215921 -5646
rect 215863 -5686 215875 -5652
rect 215863 -5692 215921 -5686
rect 215863 -5852 215921 -5846
rect 215863 -5886 215875 -5852
rect 215863 -5892 215921 -5886
rect 216050 -5901 216120 -5514
rect 216402 -5514 216436 -5513
rect 216824 -5513 216859 -5496
rect 217139 -5513 217174 -5496
rect 216824 -5514 216858 -5513
rect 216402 -5550 216472 -5514
rect 216232 -5581 216290 -5575
rect 216232 -5615 216244 -5581
rect 216419 -5584 216490 -5550
rect 216232 -5621 216290 -5615
rect 216050 -5935 216121 -5901
rect 216419 -5935 216489 -5584
rect 216601 -5652 216659 -5646
rect 216601 -5686 216613 -5652
rect 216601 -5692 216659 -5686
rect 216601 -5852 216659 -5846
rect 216601 -5886 216613 -5852
rect 216601 -5892 216659 -5886
rect 216788 -5901 216858 -5514
rect 217140 -5514 217174 -5513
rect 217562 -5513 217597 -5496
rect 217877 -5513 217912 -5496
rect 217562 -5514 217596 -5513
rect 217140 -5550 217210 -5514
rect 216970 -5581 217028 -5575
rect 216970 -5615 216982 -5581
rect 217157 -5584 217228 -5550
rect 216970 -5621 217028 -5615
rect 216788 -5935 216859 -5901
rect 217157 -5935 217227 -5584
rect 217339 -5652 217397 -5646
rect 217339 -5686 217351 -5652
rect 217339 -5692 217397 -5686
rect 217339 -5852 217397 -5846
rect 217339 -5886 217351 -5852
rect 217339 -5892 217397 -5886
rect 217526 -5901 217596 -5514
rect 217878 -5514 217912 -5513
rect 218300 -5513 218335 -5496
rect 218615 -5513 218650 -5496
rect 218300 -5514 218334 -5513
rect 217878 -5550 217948 -5514
rect 217708 -5581 217766 -5575
rect 217708 -5615 217720 -5581
rect 217895 -5584 217966 -5550
rect 217708 -5621 217766 -5615
rect 217526 -5935 217597 -5901
rect 217895 -5935 217965 -5584
rect 218077 -5652 218135 -5646
rect 218077 -5686 218089 -5652
rect 218077 -5692 218135 -5686
rect 218077 -5852 218135 -5846
rect 218077 -5886 218089 -5852
rect 218077 -5892 218135 -5886
rect 218264 -5901 218334 -5514
rect 218616 -5514 218650 -5513
rect 219038 -5513 219073 -5496
rect 219353 -5513 219388 -5496
rect 219038 -5514 219072 -5513
rect 218616 -5550 218686 -5514
rect 218446 -5581 218504 -5575
rect 218446 -5615 218458 -5581
rect 218633 -5584 218704 -5550
rect 218446 -5621 218504 -5615
rect 218264 -5935 218335 -5901
rect 218633 -5935 218703 -5584
rect 218815 -5652 218873 -5646
rect 218815 -5686 218827 -5652
rect 218815 -5692 218873 -5686
rect 218815 -5852 218873 -5846
rect 218815 -5886 218827 -5852
rect 218815 -5892 218873 -5886
rect 219002 -5901 219072 -5514
rect 219354 -5514 219388 -5513
rect 219776 -5513 219811 -5496
rect 220091 -5513 220126 -5496
rect 219776 -5514 219810 -5513
rect 219354 -5550 219424 -5514
rect 219184 -5581 219242 -5575
rect 219184 -5615 219196 -5581
rect 219371 -5584 219442 -5550
rect 219184 -5621 219242 -5615
rect 219002 -5935 219073 -5901
rect 219371 -5935 219441 -5584
rect 219553 -5652 219611 -5646
rect 219553 -5686 219565 -5652
rect 219553 -5692 219611 -5686
rect 219553 -5852 219611 -5846
rect 219553 -5886 219565 -5852
rect 219553 -5892 219611 -5886
rect 219740 -5901 219810 -5514
rect 220092 -5514 220126 -5513
rect 220514 -5513 220549 -5496
rect 220829 -5513 220864 -5496
rect 220514 -5514 220548 -5513
rect 220092 -5550 220162 -5514
rect 219922 -5581 219980 -5575
rect 219922 -5615 219934 -5581
rect 220109 -5584 220180 -5550
rect 219922 -5621 219980 -5615
rect 219740 -5935 219811 -5901
rect 220109 -5935 220179 -5584
rect 220291 -5652 220349 -5646
rect 220291 -5686 220303 -5652
rect 220291 -5692 220349 -5686
rect 220291 -5852 220349 -5846
rect 220291 -5886 220303 -5852
rect 220291 -5892 220349 -5886
rect 220478 -5901 220548 -5514
rect 220830 -5514 220864 -5513
rect 221252 -5513 221287 -5496
rect 221567 -5513 221602 -5496
rect 221252 -5514 221286 -5513
rect 220830 -5550 220900 -5514
rect 220660 -5581 220718 -5575
rect 220660 -5615 220672 -5581
rect 220847 -5584 220918 -5550
rect 220660 -5621 220718 -5615
rect 220478 -5935 220549 -5901
rect 220847 -5935 220917 -5584
rect 221029 -5652 221087 -5646
rect 221029 -5686 221041 -5652
rect 221029 -5692 221087 -5686
rect 221029 -5852 221087 -5846
rect 221029 -5886 221041 -5852
rect 221029 -5892 221087 -5886
rect 221216 -5901 221286 -5514
rect 221568 -5514 221602 -5513
rect 221990 -5513 222025 -5496
rect 222305 -5513 222340 -5496
rect 221990 -5514 222024 -5513
rect 221568 -5550 221638 -5514
rect 221398 -5581 221456 -5575
rect 221398 -5615 221410 -5581
rect 221585 -5584 221656 -5550
rect 221398 -5621 221456 -5615
rect 221216 -5935 221287 -5901
rect 221585 -5935 221655 -5584
rect 221767 -5652 221825 -5646
rect 221767 -5686 221779 -5652
rect 221767 -5692 221825 -5686
rect 221767 -5852 221825 -5846
rect 221767 -5886 221779 -5852
rect 221767 -5892 221825 -5886
rect 221954 -5901 222024 -5514
rect 222306 -5514 222340 -5513
rect 222728 -5513 222763 -5496
rect 223043 -5513 223078 -5496
rect 222728 -5514 222762 -5513
rect 222306 -5550 222376 -5514
rect 222136 -5581 222194 -5575
rect 222136 -5615 222148 -5581
rect 222323 -5584 222394 -5550
rect 222136 -5621 222194 -5615
rect 221954 -5935 222025 -5901
rect 222323 -5935 222393 -5584
rect 222505 -5652 222563 -5646
rect 222505 -5686 222517 -5652
rect 222505 -5692 222563 -5686
rect 222505 -5852 222563 -5846
rect 222505 -5886 222517 -5852
rect 222505 -5892 222563 -5886
rect 222692 -5901 222762 -5514
rect 223044 -5514 223078 -5513
rect 223466 -5513 223501 -5496
rect 223781 -5513 223816 -5496
rect 223466 -5514 223500 -5513
rect 223044 -5550 223114 -5514
rect 222874 -5581 222932 -5575
rect 222874 -5615 222886 -5581
rect 223061 -5584 223132 -5550
rect 222874 -5621 222932 -5615
rect 222692 -5935 222763 -5901
rect 223061 -5935 223131 -5584
rect 223243 -5652 223301 -5646
rect 223243 -5686 223255 -5652
rect 223243 -5692 223301 -5686
rect 223243 -5852 223301 -5846
rect 223243 -5886 223255 -5852
rect 223243 -5892 223301 -5886
rect 223430 -5901 223500 -5514
rect 223782 -5514 223816 -5513
rect 224204 -5513 224239 -5496
rect 224519 -5513 224554 -5496
rect 224204 -5514 224238 -5513
rect 223782 -5550 223852 -5514
rect 223612 -5581 223670 -5575
rect 223612 -5615 223624 -5581
rect 223799 -5584 223870 -5550
rect 223612 -5621 223670 -5615
rect 223430 -5935 223501 -5901
rect 223799 -5935 223869 -5584
rect 223981 -5652 224039 -5646
rect 223981 -5686 223993 -5652
rect 223981 -5692 224039 -5686
rect 223981 -5852 224039 -5846
rect 223981 -5886 223993 -5852
rect 223981 -5892 224039 -5886
rect 224168 -5901 224238 -5514
rect 224520 -5514 224554 -5513
rect 224942 -5513 224977 -5496
rect 225257 -5513 225292 -5496
rect 224942 -5514 224976 -5513
rect 224520 -5550 224590 -5514
rect 224350 -5581 224408 -5575
rect 224350 -5615 224362 -5581
rect 224537 -5584 224608 -5550
rect 224350 -5621 224408 -5615
rect 224168 -5935 224239 -5901
rect 224537 -5935 224607 -5584
rect 224719 -5652 224777 -5646
rect 224719 -5686 224731 -5652
rect 224719 -5692 224777 -5686
rect 224719 -5852 224777 -5846
rect 224719 -5886 224731 -5852
rect 224719 -5892 224777 -5886
rect 224906 -5901 224976 -5514
rect 225258 -5514 225292 -5513
rect 225680 -5513 225715 -5496
rect 225995 -5513 226030 -5496
rect 225680 -5514 225714 -5513
rect 225258 -5550 225328 -5514
rect 225088 -5581 225146 -5575
rect 225088 -5615 225100 -5581
rect 225275 -5584 225346 -5550
rect 225088 -5621 225146 -5615
rect 224906 -5935 224977 -5901
rect 225275 -5935 225345 -5584
rect 225457 -5652 225515 -5646
rect 225457 -5686 225469 -5652
rect 225457 -5692 225515 -5686
rect 225457 -5852 225515 -5846
rect 225457 -5886 225469 -5852
rect 225457 -5892 225515 -5886
rect 225644 -5901 225714 -5514
rect 225996 -5514 226030 -5513
rect 226418 -5513 226453 -5496
rect 226733 -5513 226768 -5496
rect 226418 -5514 226452 -5513
rect 225996 -5550 226066 -5514
rect 225826 -5581 225884 -5575
rect 225826 -5615 225838 -5581
rect 226013 -5584 226084 -5550
rect 225826 -5621 225884 -5615
rect 225644 -5935 225715 -5901
rect 226013 -5935 226083 -5584
rect 226195 -5652 226253 -5646
rect 226195 -5686 226207 -5652
rect 226195 -5692 226253 -5686
rect 226195 -5852 226253 -5846
rect 226195 -5886 226207 -5852
rect 226195 -5892 226253 -5886
rect 226382 -5901 226452 -5514
rect 226734 -5514 226768 -5513
rect 227156 -5513 227191 -5496
rect 227471 -5513 227506 -5496
rect 227156 -5514 227190 -5513
rect 226734 -5550 226804 -5514
rect 226564 -5581 226622 -5575
rect 226564 -5615 226576 -5581
rect 226751 -5584 226822 -5550
rect 226564 -5621 226622 -5615
rect 226382 -5935 226453 -5901
rect 226751 -5935 226821 -5584
rect 226933 -5652 226991 -5646
rect 226933 -5686 226945 -5652
rect 226933 -5692 226991 -5686
rect 226933 -5852 226991 -5846
rect 226933 -5886 226945 -5852
rect 226933 -5892 226991 -5886
rect 227120 -5901 227190 -5514
rect 227472 -5514 227506 -5513
rect 227894 -5513 227929 -5496
rect 228209 -5513 228244 -5496
rect 227894 -5514 227928 -5513
rect 227472 -5550 227542 -5514
rect 227302 -5581 227360 -5575
rect 227302 -5615 227314 -5581
rect 227489 -5584 227560 -5550
rect 227302 -5621 227360 -5615
rect 227120 -5935 227191 -5901
rect 227489 -5935 227559 -5584
rect 227671 -5652 227729 -5646
rect 227671 -5686 227683 -5652
rect 227671 -5692 227729 -5686
rect 227671 -5852 227729 -5846
rect 227671 -5886 227683 -5852
rect 227671 -5892 227729 -5886
rect 227858 -5901 227928 -5514
rect 228210 -5514 228244 -5513
rect 228632 -5513 228667 -5496
rect 228947 -5513 228982 -5496
rect 228632 -5514 228666 -5513
rect 228210 -5550 228280 -5514
rect 228040 -5581 228098 -5575
rect 228040 -5615 228052 -5581
rect 228227 -5584 228298 -5550
rect 228040 -5621 228098 -5615
rect 227858 -5935 227929 -5901
rect 228227 -5935 228297 -5584
rect 228409 -5652 228467 -5646
rect 228409 -5686 228421 -5652
rect 228409 -5692 228467 -5686
rect 228409 -5852 228467 -5846
rect 228409 -5886 228421 -5852
rect 228409 -5892 228467 -5886
rect 228596 -5901 228666 -5514
rect 228948 -5514 228982 -5513
rect 229370 -5513 229405 -5496
rect 229685 -5513 229720 -5496
rect 229370 -5514 229404 -5513
rect 228948 -5550 229018 -5514
rect 228778 -5581 228836 -5575
rect 228778 -5615 228790 -5581
rect 228965 -5584 229036 -5550
rect 228778 -5621 228836 -5615
rect 228596 -5935 228667 -5901
rect 228965 -5935 229035 -5584
rect 229147 -5652 229205 -5646
rect 229147 -5686 229159 -5652
rect 229147 -5692 229205 -5686
rect 229147 -5852 229205 -5846
rect 229147 -5886 229159 -5852
rect 229147 -5892 229205 -5886
rect 229334 -5901 229404 -5514
rect 229686 -5514 229720 -5513
rect 230108 -5513 230143 -5496
rect 230423 -5513 230458 -5496
rect 230108 -5514 230142 -5513
rect 229686 -5550 229756 -5514
rect 229516 -5581 229574 -5575
rect 229516 -5615 229528 -5581
rect 229703 -5584 229774 -5550
rect 229516 -5621 229574 -5615
rect 229334 -5935 229405 -5901
rect 229703 -5935 229773 -5584
rect 229885 -5652 229943 -5646
rect 229885 -5686 229897 -5652
rect 229885 -5692 229943 -5686
rect 229885 -5852 229943 -5846
rect 229885 -5886 229897 -5852
rect 229885 -5892 229943 -5886
rect 230072 -5901 230142 -5514
rect 230424 -5514 230458 -5513
rect 230846 -5513 230881 -5496
rect 231161 -5513 231196 -5496
rect 230846 -5514 230880 -5513
rect 230424 -5550 230494 -5514
rect 230254 -5581 230312 -5575
rect 230254 -5615 230266 -5581
rect 230441 -5584 230512 -5550
rect 230254 -5621 230312 -5615
rect 230072 -5935 230143 -5901
rect 230441 -5935 230511 -5584
rect 230623 -5652 230681 -5646
rect 230623 -5686 230635 -5652
rect 230623 -5692 230681 -5686
rect 230623 -5852 230681 -5846
rect 230623 -5886 230635 -5852
rect 230623 -5892 230681 -5886
rect 230810 -5901 230880 -5514
rect 231162 -5514 231196 -5513
rect 231584 -5513 231619 -5496
rect 231899 -5513 231934 -5496
rect 231584 -5514 231618 -5513
rect 231162 -5550 231232 -5514
rect 230992 -5581 231050 -5575
rect 230992 -5615 231004 -5581
rect 231179 -5584 231250 -5550
rect 230992 -5621 231050 -5615
rect 230810 -5935 230881 -5901
rect 231179 -5935 231249 -5584
rect 231361 -5652 231419 -5646
rect 231361 -5686 231373 -5652
rect 231361 -5692 231419 -5686
rect 231361 -5852 231419 -5846
rect 231361 -5886 231373 -5852
rect 231361 -5892 231419 -5886
rect 231548 -5901 231618 -5514
rect 231900 -5514 231934 -5513
rect 232322 -5513 232357 -5496
rect 232637 -5513 232672 -5496
rect 232322 -5514 232356 -5513
rect 231900 -5550 231970 -5514
rect 231730 -5581 231788 -5575
rect 231730 -5615 231742 -5581
rect 231917 -5584 231988 -5550
rect 231730 -5621 231788 -5615
rect 231548 -5935 231619 -5901
rect 231917 -5935 231987 -5584
rect 232099 -5652 232157 -5646
rect 232099 -5686 232111 -5652
rect 232099 -5692 232157 -5686
rect 232099 -5852 232157 -5846
rect 232099 -5886 232111 -5852
rect 232099 -5892 232157 -5886
rect 232286 -5901 232356 -5514
rect 232638 -5514 232672 -5513
rect 233060 -5513 233095 -5496
rect 233375 -5513 233410 -5496
rect 233060 -5514 233094 -5513
rect 232638 -5550 232708 -5514
rect 232468 -5581 232526 -5575
rect 232468 -5615 232480 -5581
rect 232655 -5584 232726 -5550
rect 232468 -5621 232526 -5615
rect 232286 -5935 232357 -5901
rect 232655 -5935 232725 -5584
rect 232837 -5652 232895 -5646
rect 232837 -5686 232849 -5652
rect 232837 -5692 232895 -5686
rect 232837 -5852 232895 -5846
rect 232837 -5886 232849 -5852
rect 232837 -5892 232895 -5886
rect 233024 -5901 233094 -5514
rect 233376 -5514 233410 -5513
rect 233798 -5513 233833 -5496
rect 234113 -5513 234148 -5496
rect 233798 -5514 233832 -5513
rect 233376 -5550 233446 -5514
rect 233206 -5581 233264 -5575
rect 233206 -5615 233218 -5581
rect 233393 -5584 233464 -5550
rect 233206 -5621 233264 -5615
rect 233024 -5935 233095 -5901
rect 233393 -5935 233463 -5584
rect 233575 -5652 233633 -5646
rect 233575 -5686 233587 -5652
rect 233575 -5692 233633 -5686
rect 233575 -5852 233633 -5846
rect 233575 -5886 233587 -5852
rect 233575 -5892 233633 -5886
rect 233762 -5901 233832 -5514
rect 234114 -5514 234148 -5513
rect 234536 -5513 234571 -5496
rect 234851 -5513 234886 -5496
rect 234536 -5514 234570 -5513
rect 234114 -5550 234184 -5514
rect 233944 -5581 234002 -5575
rect 233944 -5615 233956 -5581
rect 234131 -5584 234202 -5550
rect 233944 -5621 234002 -5615
rect 233762 -5935 233833 -5901
rect 234131 -5935 234201 -5584
rect 234313 -5652 234371 -5646
rect 234313 -5686 234325 -5652
rect 234313 -5692 234371 -5686
rect 234313 -5852 234371 -5846
rect 234313 -5886 234325 -5852
rect 234313 -5892 234371 -5886
rect 234500 -5901 234570 -5514
rect 234852 -5514 234886 -5513
rect 235274 -5513 235309 -5496
rect 235589 -5513 235624 -5496
rect 235274 -5514 235308 -5513
rect 234852 -5550 234922 -5514
rect 234682 -5581 234740 -5575
rect 234682 -5615 234694 -5581
rect 234869 -5584 234940 -5550
rect 234682 -5621 234740 -5615
rect 234500 -5935 234571 -5901
rect 234869 -5935 234939 -5584
rect 235051 -5652 235109 -5646
rect 235051 -5686 235063 -5652
rect 235051 -5692 235109 -5686
rect 235051 -5852 235109 -5846
rect 235051 -5886 235063 -5852
rect 235051 -5892 235109 -5886
rect 235238 -5901 235308 -5514
rect 235590 -5514 235624 -5513
rect 236012 -5513 236047 -5496
rect 236327 -5513 236362 -5496
rect 236012 -5514 236046 -5513
rect 235590 -5550 235660 -5514
rect 235420 -5581 235478 -5575
rect 235420 -5615 235432 -5581
rect 235607 -5584 235678 -5550
rect 235420 -5621 235478 -5615
rect 235238 -5935 235309 -5901
rect 235607 -5935 235677 -5584
rect 235789 -5652 235847 -5646
rect 235789 -5686 235801 -5652
rect 235789 -5692 235847 -5686
rect 235789 -5852 235847 -5846
rect 235789 -5886 235801 -5852
rect 235789 -5892 235847 -5886
rect 235976 -5901 236046 -5514
rect 236328 -5514 236362 -5513
rect 236750 -5513 236785 -5496
rect 237065 -5513 237100 -5496
rect 236750 -5514 236784 -5513
rect 236328 -5550 236398 -5514
rect 236158 -5581 236216 -5575
rect 236158 -5615 236170 -5581
rect 236345 -5584 236416 -5550
rect 236158 -5621 236216 -5615
rect 235976 -5935 236047 -5901
rect 236345 -5935 236415 -5584
rect 236527 -5652 236585 -5646
rect 236527 -5686 236539 -5652
rect 236527 -5692 236585 -5686
rect 236527 -5852 236585 -5846
rect 236527 -5886 236539 -5852
rect 236527 -5892 236585 -5886
rect 236714 -5901 236784 -5514
rect 237066 -5514 237100 -5513
rect 237488 -5513 237523 -5496
rect 237803 -5513 237838 -5496
rect 237488 -5514 237522 -5513
rect 237066 -5550 237136 -5514
rect 236896 -5581 236954 -5575
rect 236896 -5615 236908 -5581
rect 237083 -5584 237154 -5550
rect 236896 -5621 236954 -5615
rect 236714 -5935 236785 -5901
rect 237083 -5935 237153 -5584
rect 237265 -5652 237323 -5646
rect 237265 -5686 237277 -5652
rect 237265 -5692 237323 -5686
rect 237265 -5852 237323 -5846
rect 237265 -5886 237277 -5852
rect 237265 -5892 237323 -5886
rect 237452 -5901 237522 -5514
rect 237804 -5514 237838 -5513
rect 238226 -5513 238261 -5496
rect 238541 -5513 238576 -5496
rect 238226 -5514 238260 -5513
rect 237804 -5550 237874 -5514
rect 237634 -5581 237692 -5575
rect 237634 -5615 237646 -5581
rect 237821 -5584 237892 -5550
rect 237634 -5621 237692 -5615
rect 237452 -5935 237523 -5901
rect 237821 -5935 237891 -5584
rect 238003 -5652 238061 -5646
rect 238003 -5686 238015 -5652
rect 238003 -5692 238061 -5686
rect 238003 -5852 238061 -5846
rect 238003 -5886 238015 -5852
rect 238003 -5892 238061 -5886
rect 238190 -5901 238260 -5514
rect 238542 -5514 238576 -5513
rect 238964 -5513 238999 -5496
rect 239279 -5513 239314 -5496
rect 238964 -5514 238998 -5513
rect 238542 -5550 238612 -5514
rect 238372 -5581 238430 -5575
rect 238372 -5615 238384 -5581
rect 238559 -5584 238630 -5550
rect 238372 -5621 238430 -5615
rect 238190 -5935 238261 -5901
rect 238559 -5935 238629 -5584
rect 238741 -5652 238799 -5646
rect 238741 -5686 238753 -5652
rect 238741 -5692 238799 -5686
rect 238741 -5852 238799 -5846
rect 238741 -5886 238753 -5852
rect 238741 -5892 238799 -5886
rect 238928 -5901 238998 -5514
rect 239280 -5514 239314 -5513
rect 239702 -5513 239737 -5496
rect 240017 -5513 240052 -5496
rect 239702 -5514 239736 -5513
rect 239280 -5550 239350 -5514
rect 239110 -5581 239168 -5575
rect 239110 -5615 239122 -5581
rect 239297 -5584 239368 -5550
rect 239110 -5621 239168 -5615
rect 238928 -5935 238999 -5901
rect 239297 -5935 239367 -5584
rect 239479 -5652 239537 -5646
rect 239479 -5686 239491 -5652
rect 239479 -5692 239537 -5686
rect 239479 -5852 239537 -5846
rect 239479 -5886 239491 -5852
rect 239479 -5892 239537 -5886
rect 239666 -5901 239736 -5514
rect 240018 -5514 240052 -5513
rect 240440 -5513 240475 -5496
rect 240755 -5513 240790 -5496
rect 240440 -5514 240474 -5513
rect 240018 -5550 240088 -5514
rect 239848 -5581 239906 -5575
rect 239848 -5615 239860 -5581
rect 240035 -5584 240106 -5550
rect 239848 -5621 239906 -5615
rect 239666 -5935 239737 -5901
rect 240035 -5935 240105 -5584
rect 240217 -5652 240275 -5646
rect 240217 -5686 240229 -5652
rect 240217 -5692 240275 -5686
rect 240217 -5852 240275 -5846
rect 240217 -5886 240229 -5852
rect 240217 -5892 240275 -5886
rect 240404 -5901 240474 -5514
rect 240756 -5514 240790 -5513
rect 241178 -5513 241213 -5496
rect 241493 -5513 241528 -5496
rect 241178 -5514 241212 -5513
rect 240756 -5550 240826 -5514
rect 240586 -5581 240644 -5575
rect 240586 -5615 240598 -5581
rect 240773 -5584 240844 -5550
rect 240586 -5621 240644 -5615
rect 240404 -5935 240475 -5901
rect 240773 -5935 240843 -5584
rect 240955 -5652 241013 -5646
rect 240955 -5686 240967 -5652
rect 240955 -5692 241013 -5686
rect 240955 -5852 241013 -5846
rect 240955 -5886 240967 -5852
rect 240955 -5892 241013 -5886
rect 241142 -5901 241212 -5514
rect 241494 -5514 241528 -5513
rect 241916 -5513 241951 -5496
rect 242231 -5513 242266 -5496
rect 241916 -5514 241950 -5513
rect 241494 -5550 241564 -5514
rect 241324 -5581 241382 -5575
rect 241324 -5615 241336 -5581
rect 241511 -5584 241582 -5550
rect 241324 -5621 241382 -5615
rect 241142 -5935 241213 -5901
rect 241511 -5935 241581 -5584
rect 241693 -5652 241751 -5646
rect 241693 -5686 241705 -5652
rect 241693 -5692 241751 -5686
rect 241693 -5852 241751 -5846
rect 241693 -5886 241705 -5852
rect 241693 -5892 241751 -5886
rect 241880 -5901 241950 -5514
rect 242232 -5514 242266 -5513
rect 242654 -5513 242689 -5496
rect 242969 -5513 243004 -5496
rect 242654 -5514 242688 -5513
rect 242232 -5550 242302 -5514
rect 242062 -5581 242120 -5575
rect 242062 -5615 242074 -5581
rect 242249 -5584 242320 -5550
rect 242062 -5621 242120 -5615
rect 241880 -5935 241951 -5901
rect 242249 -5935 242319 -5584
rect 242431 -5652 242489 -5646
rect 242431 -5686 242443 -5652
rect 242431 -5692 242489 -5686
rect 242431 -5852 242489 -5846
rect 242431 -5886 242443 -5852
rect 242431 -5892 242489 -5886
rect 242618 -5901 242688 -5514
rect 242970 -5514 243004 -5513
rect 243392 -5513 243427 -5496
rect 243707 -5513 243742 -5496
rect 243392 -5514 243426 -5513
rect 242970 -5550 243040 -5514
rect 242800 -5581 242858 -5575
rect 242800 -5615 242812 -5581
rect 242987 -5584 243058 -5550
rect 242800 -5621 242858 -5615
rect 242618 -5935 242689 -5901
rect 242987 -5935 243057 -5584
rect 243169 -5652 243227 -5646
rect 243169 -5686 243181 -5652
rect 243169 -5692 243227 -5686
rect 243169 -5852 243227 -5846
rect 243169 -5886 243181 -5852
rect 243169 -5892 243227 -5886
rect 243356 -5901 243426 -5514
rect 243708 -5514 243742 -5513
rect 244130 -5513 244165 -5496
rect 244445 -5513 244480 -5496
rect 244130 -5514 244164 -5513
rect 243708 -5550 243778 -5514
rect 243538 -5581 243596 -5575
rect 243538 -5615 243550 -5581
rect 243725 -5584 243796 -5550
rect 243538 -5621 243596 -5615
rect 243356 -5935 243427 -5901
rect 243725 -5935 243795 -5584
rect 243907 -5652 243965 -5646
rect 243907 -5686 243919 -5652
rect 243907 -5692 243965 -5686
rect 243907 -5852 243965 -5846
rect 243907 -5886 243919 -5852
rect 243907 -5892 243965 -5886
rect 244094 -5901 244164 -5514
rect 244446 -5514 244480 -5513
rect 244868 -5513 244903 -5496
rect 245183 -5513 245218 -5496
rect 244868 -5514 244902 -5513
rect 244446 -5550 244516 -5514
rect 244276 -5581 244334 -5575
rect 244276 -5615 244288 -5581
rect 244463 -5584 244534 -5550
rect 244276 -5621 244334 -5615
rect 244094 -5935 244165 -5901
rect 244463 -5935 244533 -5584
rect 244645 -5652 244703 -5646
rect 244645 -5686 244657 -5652
rect 244645 -5692 244703 -5686
rect 244645 -5852 244703 -5846
rect 244645 -5886 244657 -5852
rect 244645 -5892 244703 -5886
rect 244832 -5901 244902 -5514
rect 245184 -5514 245218 -5513
rect 245606 -5513 245641 -5496
rect 245921 -5513 245956 -5496
rect 245606 -5514 245640 -5513
rect 245184 -5550 245254 -5514
rect 245014 -5581 245072 -5575
rect 245014 -5615 245026 -5581
rect 245201 -5584 245272 -5550
rect 245014 -5621 245072 -5615
rect 244832 -5935 244903 -5901
rect 245201 -5935 245271 -5584
rect 245383 -5652 245441 -5646
rect 245383 -5686 245395 -5652
rect 245383 -5692 245441 -5686
rect 245383 -5852 245441 -5846
rect 245383 -5886 245395 -5852
rect 245383 -5892 245441 -5886
rect 245570 -5901 245640 -5514
rect 245922 -5514 245956 -5513
rect 246344 -5513 246379 -5496
rect 246659 -5513 246694 -5496
rect 246344 -5514 246378 -5513
rect 245922 -5550 245992 -5514
rect 245752 -5581 245810 -5575
rect 245752 -5615 245764 -5581
rect 245939 -5584 246010 -5550
rect 245752 -5621 245810 -5615
rect 245570 -5935 245641 -5901
rect 245939 -5935 246009 -5584
rect 246121 -5652 246179 -5646
rect 246121 -5686 246133 -5652
rect 246121 -5692 246179 -5686
rect 246121 -5852 246179 -5846
rect 246121 -5886 246133 -5852
rect 246121 -5892 246179 -5886
rect 246308 -5901 246378 -5514
rect 246660 -5514 246694 -5513
rect 247082 -5513 247117 -5496
rect 247397 -5513 247432 -5496
rect 247082 -5514 247116 -5513
rect 246660 -5550 246730 -5514
rect 246490 -5581 246548 -5575
rect 246490 -5615 246502 -5581
rect 246677 -5584 246748 -5550
rect 246490 -5621 246548 -5615
rect 246308 -5935 246379 -5901
rect 246677 -5935 246747 -5584
rect 246859 -5652 246917 -5646
rect 246859 -5686 246871 -5652
rect 246859 -5692 246917 -5686
rect 246859 -5852 246917 -5846
rect 246859 -5886 246871 -5852
rect 246859 -5892 246917 -5886
rect 247046 -5901 247116 -5514
rect 247398 -5514 247432 -5513
rect 247820 -5513 247855 -5496
rect 248135 -5513 248170 -5496
rect 247820 -5514 247854 -5513
rect 247398 -5550 247468 -5514
rect 247228 -5581 247286 -5575
rect 247228 -5615 247240 -5581
rect 247415 -5584 247486 -5550
rect 247228 -5621 247286 -5615
rect 247046 -5935 247117 -5901
rect 247415 -5935 247485 -5584
rect 247597 -5652 247655 -5646
rect 247597 -5686 247609 -5652
rect 247597 -5692 247655 -5686
rect 247597 -5852 247655 -5846
rect 247597 -5886 247609 -5852
rect 247597 -5892 247655 -5886
rect 247784 -5901 247854 -5514
rect 248136 -5514 248170 -5513
rect 248558 -5513 248593 -5496
rect 248873 -5513 248908 -5496
rect 248558 -5514 248592 -5513
rect 248136 -5550 248206 -5514
rect 247966 -5581 248024 -5575
rect 247966 -5615 247978 -5581
rect 248153 -5584 248224 -5550
rect 247966 -5621 248024 -5615
rect 247784 -5935 247855 -5901
rect 248153 -5935 248223 -5584
rect 248335 -5652 248393 -5646
rect 248335 -5686 248347 -5652
rect 248335 -5692 248393 -5686
rect 248335 -5852 248393 -5846
rect 248335 -5886 248347 -5852
rect 248335 -5892 248393 -5886
rect 248522 -5901 248592 -5514
rect 248874 -5514 248908 -5513
rect 249296 -5513 249331 -5496
rect 249611 -5513 249646 -5496
rect 249296 -5514 249330 -5513
rect 248874 -5550 248944 -5514
rect 248704 -5581 248762 -5575
rect 248704 -5615 248716 -5581
rect 248891 -5584 248962 -5550
rect 248704 -5621 248762 -5615
rect 248522 -5935 248593 -5901
rect 248891 -5935 248961 -5584
rect 249073 -5652 249131 -5646
rect 249073 -5686 249085 -5652
rect 249073 -5692 249131 -5686
rect 249073 -5852 249131 -5846
rect 249073 -5886 249085 -5852
rect 249073 -5892 249131 -5886
rect 249260 -5901 249330 -5514
rect 249612 -5514 249646 -5513
rect 250034 -5513 250069 -5496
rect 250349 -5513 250384 -5496
rect 250034 -5514 250068 -5513
rect 249612 -5550 249682 -5514
rect 249442 -5581 249500 -5575
rect 249442 -5615 249454 -5581
rect 249629 -5584 249700 -5550
rect 249442 -5621 249500 -5615
rect 249260 -5935 249331 -5901
rect 249629 -5935 249699 -5584
rect 249811 -5652 249869 -5646
rect 249811 -5686 249823 -5652
rect 249811 -5692 249869 -5686
rect 249811 -5852 249869 -5846
rect 249811 -5886 249823 -5852
rect 249811 -5892 249869 -5886
rect 249998 -5901 250068 -5514
rect 250350 -5514 250384 -5513
rect 250772 -5513 250807 -5496
rect 251087 -5513 251122 -5496
rect 250772 -5514 250806 -5513
rect 250350 -5550 250420 -5514
rect 250180 -5581 250238 -5575
rect 250180 -5615 250192 -5581
rect 250367 -5584 250438 -5550
rect 250180 -5621 250238 -5615
rect 249998 -5935 250069 -5901
rect 250367 -5935 250437 -5584
rect 250549 -5652 250607 -5646
rect 250549 -5686 250561 -5652
rect 250549 -5692 250607 -5686
rect 250549 -5852 250607 -5846
rect 250549 -5886 250561 -5852
rect 250549 -5892 250607 -5886
rect 250736 -5901 250806 -5514
rect 251088 -5514 251122 -5513
rect 251510 -5513 251545 -5496
rect 251825 -5513 251860 -5496
rect 251510 -5514 251544 -5513
rect 251088 -5550 251158 -5514
rect 250918 -5581 250976 -5575
rect 250918 -5615 250930 -5581
rect 251105 -5584 251176 -5550
rect 250918 -5621 250976 -5615
rect 250736 -5935 250807 -5901
rect 251105 -5935 251175 -5584
rect 251287 -5652 251345 -5646
rect 251287 -5686 251299 -5652
rect 251287 -5692 251345 -5686
rect 251287 -5852 251345 -5846
rect 251287 -5886 251299 -5852
rect 251287 -5892 251345 -5886
rect 251474 -5901 251544 -5514
rect 251826 -5514 251860 -5513
rect 252248 -5513 252283 -5496
rect 252563 -5513 252598 -5496
rect 252248 -5514 252282 -5513
rect 251826 -5550 251896 -5514
rect 251656 -5581 251714 -5575
rect 251656 -5615 251668 -5581
rect 251843 -5584 251914 -5550
rect 251656 -5621 251714 -5615
rect 251474 -5935 251545 -5901
rect 251843 -5935 251913 -5584
rect 252025 -5652 252083 -5646
rect 252025 -5686 252037 -5652
rect 252025 -5692 252083 -5686
rect 252025 -5852 252083 -5846
rect 252025 -5886 252037 -5852
rect 252025 -5892 252083 -5886
rect 252212 -5901 252282 -5514
rect 252564 -5514 252598 -5513
rect 252986 -5513 253021 -5496
rect 253301 -5513 253336 -5496
rect 252986 -5514 253020 -5513
rect 252564 -5550 252634 -5514
rect 252394 -5581 252452 -5575
rect 252394 -5615 252406 -5581
rect 252581 -5584 252652 -5550
rect 252394 -5621 252452 -5615
rect 252212 -5935 252283 -5901
rect 252581 -5935 252651 -5584
rect 252763 -5652 252821 -5646
rect 252763 -5686 252775 -5652
rect 252763 -5692 252821 -5686
rect 252763 -5852 252821 -5846
rect 252763 -5886 252775 -5852
rect 252763 -5892 252821 -5886
rect 252950 -5901 253020 -5514
rect 253302 -5514 253336 -5513
rect 253724 -5513 253759 -5496
rect 254039 -5513 254074 -5496
rect 253724 -5514 253758 -5513
rect 253302 -5550 253372 -5514
rect 253132 -5581 253190 -5575
rect 253132 -5615 253144 -5581
rect 253319 -5584 253390 -5550
rect 253132 -5621 253190 -5615
rect 252950 -5935 253021 -5901
rect 253319 -5935 253389 -5584
rect 253501 -5652 253559 -5646
rect 253501 -5686 253513 -5652
rect 253501 -5692 253559 -5686
rect 253501 -5852 253559 -5846
rect 253501 -5886 253513 -5852
rect 253501 -5892 253559 -5886
rect 253688 -5901 253758 -5514
rect 254040 -5514 254074 -5513
rect 254462 -5513 254497 -5496
rect 254777 -5513 254812 -5496
rect 254462 -5514 254496 -5513
rect 254040 -5550 254110 -5514
rect 253870 -5581 253928 -5575
rect 253870 -5615 253882 -5581
rect 254057 -5584 254128 -5550
rect 253870 -5621 253928 -5615
rect 253688 -5935 253759 -5901
rect 254057 -5935 254127 -5584
rect 254239 -5652 254297 -5646
rect 254239 -5686 254251 -5652
rect 254239 -5692 254297 -5686
rect 254239 -5852 254297 -5846
rect 254239 -5886 254251 -5852
rect 254239 -5892 254297 -5886
rect 254426 -5901 254496 -5514
rect 254778 -5514 254812 -5513
rect 255200 -5513 255235 -5496
rect 255515 -5513 255550 -5496
rect 255200 -5514 255234 -5513
rect 254778 -5550 254848 -5514
rect 254608 -5581 254666 -5575
rect 254608 -5615 254620 -5581
rect 254795 -5584 254866 -5550
rect 254608 -5621 254666 -5615
rect 254426 -5935 254497 -5901
rect 254795 -5935 254865 -5584
rect 254977 -5652 255035 -5646
rect 254977 -5686 254989 -5652
rect 254977 -5692 255035 -5686
rect 254977 -5852 255035 -5846
rect 254977 -5886 254989 -5852
rect 254977 -5892 255035 -5886
rect 255164 -5901 255234 -5514
rect 255516 -5514 255550 -5513
rect 255938 -5513 255973 -5496
rect 256253 -5513 256288 -5496
rect 255938 -5514 255972 -5513
rect 255516 -5550 255586 -5514
rect 255346 -5581 255404 -5575
rect 255346 -5615 255358 -5581
rect 255533 -5584 255604 -5550
rect 255346 -5621 255404 -5615
rect 255164 -5935 255235 -5901
rect 255533 -5935 255603 -5584
rect 255715 -5652 255773 -5646
rect 255715 -5686 255727 -5652
rect 255715 -5692 255773 -5686
rect 255715 -5852 255773 -5846
rect 255715 -5886 255727 -5852
rect 255715 -5892 255773 -5886
rect 255902 -5901 255972 -5514
rect 256254 -5514 256288 -5513
rect 256676 -5513 256711 -5496
rect 256991 -5513 257026 -5496
rect 256676 -5514 256710 -5513
rect 256254 -5550 256324 -5514
rect 256084 -5581 256142 -5575
rect 256084 -5615 256096 -5581
rect 256271 -5584 256342 -5550
rect 256084 -5621 256142 -5615
rect 255902 -5935 255973 -5901
rect 256271 -5935 256341 -5584
rect 256453 -5652 256511 -5646
rect 256453 -5686 256465 -5652
rect 256453 -5692 256511 -5686
rect 256453 -5852 256511 -5846
rect 256453 -5886 256465 -5852
rect 256453 -5892 256511 -5886
rect 256640 -5901 256710 -5514
rect 256992 -5514 257026 -5513
rect 257414 -5513 257449 -5496
rect 257729 -5513 257764 -5496
rect 257414 -5514 257448 -5513
rect 256992 -5550 257062 -5514
rect 256822 -5581 256880 -5575
rect 256822 -5615 256834 -5581
rect 257009 -5584 257080 -5550
rect 256822 -5621 256880 -5615
rect 256640 -5935 256711 -5901
rect 257009 -5935 257079 -5584
rect 257191 -5652 257249 -5646
rect 257191 -5686 257203 -5652
rect 257191 -5692 257249 -5686
rect 257191 -5852 257249 -5846
rect 257191 -5886 257203 -5852
rect 257191 -5892 257249 -5886
rect 257378 -5901 257448 -5514
rect 257730 -5514 257764 -5513
rect 258152 -5513 258187 -5496
rect 258467 -5513 258502 -5496
rect 258152 -5514 258186 -5513
rect 257730 -5550 257800 -5514
rect 257560 -5581 257618 -5575
rect 257560 -5615 257572 -5581
rect 257747 -5584 257818 -5550
rect 257560 -5621 257618 -5615
rect 257378 -5935 257449 -5901
rect 257747 -5935 257817 -5584
rect 257929 -5652 257987 -5646
rect 257929 -5686 257941 -5652
rect 257929 -5692 257987 -5686
rect 257929 -5852 257987 -5846
rect 257929 -5886 257941 -5852
rect 257929 -5892 257987 -5886
rect 258116 -5901 258186 -5514
rect 258468 -5514 258502 -5513
rect 258890 -5513 258925 -5496
rect 259205 -5513 259240 -5496
rect 258890 -5514 258924 -5513
rect 258468 -5550 258538 -5514
rect 258298 -5581 258356 -5575
rect 258298 -5615 258310 -5581
rect 258485 -5584 258556 -5550
rect 258298 -5621 258356 -5615
rect 258116 -5935 258187 -5901
rect 258485 -5935 258555 -5584
rect 258667 -5652 258725 -5646
rect 258667 -5686 258679 -5652
rect 258667 -5692 258725 -5686
rect 258667 -5852 258725 -5846
rect 258667 -5886 258679 -5852
rect 258667 -5892 258725 -5886
rect 258854 -5901 258924 -5514
rect 259206 -5514 259240 -5513
rect 259628 -5513 259663 -5496
rect 259943 -5513 259978 -5496
rect 259628 -5514 259662 -5513
rect 259206 -5550 259276 -5514
rect 259036 -5581 259094 -5575
rect 259036 -5615 259048 -5581
rect 259223 -5584 259294 -5550
rect 259036 -5621 259094 -5615
rect 258854 -5935 258925 -5901
rect 259223 -5935 259293 -5584
rect 259405 -5652 259463 -5646
rect 259405 -5686 259417 -5652
rect 259405 -5692 259463 -5686
rect 259405 -5852 259463 -5846
rect 259405 -5886 259417 -5852
rect 259405 -5892 259463 -5886
rect 259592 -5901 259662 -5514
rect 259944 -5514 259978 -5513
rect 260366 -5513 260401 -5496
rect 260681 -5513 260716 -5496
rect 260366 -5514 260400 -5513
rect 259944 -5550 260014 -5514
rect 259774 -5581 259832 -5575
rect 259774 -5615 259786 -5581
rect 259961 -5584 260032 -5550
rect 259774 -5621 259832 -5615
rect 259592 -5935 259663 -5901
rect 259961 -5935 260031 -5584
rect 260143 -5652 260201 -5646
rect 260143 -5686 260155 -5652
rect 260143 -5692 260201 -5686
rect 260143 -5852 260201 -5846
rect 260143 -5886 260155 -5852
rect 260143 -5892 260201 -5886
rect 260330 -5901 260400 -5514
rect 260682 -5514 260716 -5513
rect 261104 -5513 261139 -5496
rect 261419 -5513 261454 -5496
rect 261104 -5514 261138 -5513
rect 260682 -5550 260752 -5514
rect 260512 -5581 260570 -5575
rect 260512 -5615 260524 -5581
rect 260699 -5584 260770 -5550
rect 260512 -5621 260570 -5615
rect 260330 -5935 260401 -5901
rect 260699 -5935 260769 -5584
rect 260881 -5652 260939 -5646
rect 260881 -5686 260893 -5652
rect 260881 -5692 260939 -5686
rect 260881 -5852 260939 -5846
rect 260881 -5886 260893 -5852
rect 260881 -5892 260939 -5886
rect 261068 -5901 261138 -5514
rect 261420 -5514 261454 -5513
rect 261842 -5513 261877 -5496
rect 262157 -5513 262192 -5496
rect 261842 -5514 261876 -5513
rect 261420 -5550 261490 -5514
rect 261250 -5581 261308 -5575
rect 261250 -5615 261262 -5581
rect 261437 -5584 261508 -5550
rect 261250 -5621 261308 -5615
rect 261068 -5935 261139 -5901
rect 261437 -5935 261507 -5584
rect 261619 -5652 261677 -5646
rect 261619 -5686 261631 -5652
rect 261619 -5692 261677 -5686
rect 261619 -5852 261677 -5846
rect 261619 -5886 261631 -5852
rect 261619 -5892 261677 -5886
rect 261806 -5901 261876 -5514
rect 262158 -5514 262192 -5513
rect 262580 -5513 262615 -5496
rect 262895 -5513 262930 -5496
rect 262580 -5514 262614 -5513
rect 262158 -5550 262228 -5514
rect 261988 -5581 262046 -5575
rect 261988 -5615 262000 -5581
rect 262175 -5584 262246 -5550
rect 261988 -5621 262046 -5615
rect 261806 -5935 261877 -5901
rect 262175 -5935 262245 -5584
rect 262357 -5652 262415 -5646
rect 262357 -5686 262369 -5652
rect 262357 -5692 262415 -5686
rect 262357 -5852 262415 -5846
rect 262357 -5886 262369 -5852
rect 262357 -5892 262415 -5886
rect 262544 -5901 262614 -5514
rect 262896 -5514 262930 -5513
rect 263318 -5513 263353 -5496
rect 263633 -5513 263668 -5496
rect 263318 -5514 263352 -5513
rect 262896 -5550 262966 -5514
rect 262726 -5581 262784 -5575
rect 262726 -5615 262738 -5581
rect 262913 -5584 262984 -5550
rect 262726 -5621 262784 -5615
rect 262544 -5935 262615 -5901
rect 262913 -5935 262983 -5584
rect 263095 -5652 263153 -5646
rect 263095 -5686 263107 -5652
rect 263095 -5692 263153 -5686
rect 263095 -5852 263153 -5846
rect 263095 -5886 263107 -5852
rect 263095 -5892 263153 -5886
rect 263282 -5901 263352 -5514
rect 263634 -5514 263668 -5513
rect 264056 -5513 264091 -5496
rect 264371 -5513 264406 -5496
rect 264056 -5514 264090 -5513
rect 263634 -5550 263704 -5514
rect 263464 -5581 263522 -5575
rect 263464 -5615 263476 -5581
rect 263651 -5584 263722 -5550
rect 263464 -5621 263522 -5615
rect 263282 -5935 263353 -5901
rect 263651 -5935 263721 -5584
rect 263833 -5652 263891 -5646
rect 263833 -5686 263845 -5652
rect 263833 -5692 263891 -5686
rect 263833 -5852 263891 -5846
rect 263833 -5886 263845 -5852
rect 263833 -5892 263891 -5886
rect 264020 -5901 264090 -5514
rect 264372 -5514 264406 -5513
rect 264794 -5513 264829 -5496
rect 265109 -5513 265144 -5496
rect 264794 -5514 264828 -5513
rect 264372 -5550 264442 -5514
rect 264202 -5581 264260 -5575
rect 264202 -5615 264214 -5581
rect 264389 -5584 264460 -5550
rect 264202 -5621 264260 -5615
rect 264020 -5935 264091 -5901
rect 264389 -5935 264459 -5584
rect 264571 -5652 264629 -5646
rect 264571 -5686 264583 -5652
rect 264571 -5692 264629 -5686
rect 264571 -5852 264629 -5846
rect 264571 -5886 264583 -5852
rect 264571 -5892 264629 -5886
rect 264758 -5901 264828 -5514
rect 265110 -5514 265144 -5513
rect 265532 -5513 265567 -5496
rect 265847 -5513 265882 -5496
rect 265532 -5514 265566 -5513
rect 265110 -5550 265180 -5514
rect 264940 -5581 264998 -5575
rect 264940 -5615 264952 -5581
rect 265127 -5584 265198 -5550
rect 264940 -5621 264998 -5615
rect 264758 -5935 264829 -5901
rect 265127 -5935 265197 -5584
rect 265309 -5652 265367 -5646
rect 265309 -5686 265321 -5652
rect 265309 -5692 265367 -5686
rect 265309 -5852 265367 -5846
rect 265309 -5886 265321 -5852
rect 265309 -5892 265367 -5886
rect 265496 -5901 265566 -5514
rect 265848 -5514 265882 -5513
rect 266270 -5513 266305 -5496
rect 266585 -5513 266620 -5496
rect 266270 -5514 266304 -5513
rect 265848 -5550 265918 -5514
rect 265678 -5581 265736 -5575
rect 265678 -5615 265690 -5581
rect 265865 -5584 265936 -5550
rect 265678 -5621 265736 -5615
rect 265496 -5935 265567 -5901
rect 265865 -5935 265935 -5584
rect 266047 -5652 266105 -5646
rect 266047 -5686 266059 -5652
rect 266047 -5692 266105 -5686
rect 266047 -5852 266105 -5846
rect 266047 -5886 266059 -5852
rect 266047 -5892 266105 -5886
rect 266234 -5901 266304 -5514
rect 266586 -5514 266620 -5513
rect 267008 -5513 267043 -5496
rect 267323 -5513 267358 -5496
rect 267008 -5514 267042 -5513
rect 266586 -5550 266656 -5514
rect 266416 -5581 266474 -5575
rect 266416 -5615 266428 -5581
rect 266603 -5584 266674 -5550
rect 266416 -5621 266474 -5615
rect 266234 -5935 266305 -5901
rect 266603 -5935 266673 -5584
rect 266785 -5652 266843 -5646
rect 266785 -5686 266797 -5652
rect 266785 -5692 266843 -5686
rect 266785 -5852 266843 -5846
rect 266785 -5886 266797 -5852
rect 266785 -5892 266843 -5886
rect 266972 -5901 267042 -5514
rect 267324 -5514 267358 -5513
rect 267746 -5513 267781 -5496
rect 268061 -5513 268096 -5496
rect 267746 -5514 267780 -5513
rect 267324 -5550 267394 -5514
rect 267154 -5581 267212 -5575
rect 267154 -5615 267166 -5581
rect 267341 -5584 267412 -5550
rect 267154 -5621 267212 -5615
rect 266972 -5935 267043 -5901
rect 267341 -5935 267411 -5584
rect 267523 -5652 267581 -5646
rect 267523 -5686 267535 -5652
rect 267523 -5692 267581 -5686
rect 267523 -5852 267581 -5846
rect 267523 -5886 267535 -5852
rect 267523 -5892 267581 -5886
rect 267710 -5901 267780 -5514
rect 268062 -5514 268096 -5513
rect 268484 -5513 268519 -5496
rect 268799 -5513 268834 -5496
rect 268484 -5514 268518 -5513
rect 268062 -5550 268132 -5514
rect 267892 -5581 267950 -5575
rect 267892 -5615 267904 -5581
rect 268079 -5584 268150 -5550
rect 267892 -5621 267950 -5615
rect 267710 -5935 267781 -5901
rect 268079 -5935 268149 -5584
rect 268261 -5652 268319 -5646
rect 268261 -5686 268273 -5652
rect 268261 -5692 268319 -5686
rect 268261 -5852 268319 -5846
rect 268261 -5886 268273 -5852
rect 268261 -5892 268319 -5886
rect 268448 -5901 268518 -5514
rect 268800 -5514 268834 -5513
rect 269222 -5513 269257 -5496
rect 269537 -5513 269572 -5496
rect 269222 -5514 269256 -5513
rect 268800 -5550 268870 -5514
rect 268630 -5581 268688 -5575
rect 268630 -5615 268642 -5581
rect 268817 -5584 268888 -5550
rect 268630 -5621 268688 -5615
rect 268448 -5935 268519 -5901
rect 268817 -5935 268887 -5584
rect 268999 -5652 269057 -5646
rect 268999 -5686 269011 -5652
rect 268999 -5692 269057 -5686
rect 268999 -5852 269057 -5846
rect 268999 -5886 269011 -5852
rect 268999 -5892 269057 -5886
rect 269186 -5901 269256 -5514
rect 269538 -5514 269572 -5513
rect 269960 -5513 269995 -5496
rect 270275 -5513 270310 -5496
rect 269960 -5514 269994 -5513
rect 269538 -5550 269608 -5514
rect 269368 -5581 269426 -5575
rect 269368 -5615 269380 -5581
rect 269555 -5584 269626 -5550
rect 269368 -5621 269426 -5615
rect 269186 -5935 269257 -5901
rect 269555 -5935 269625 -5584
rect 269737 -5652 269795 -5646
rect 269737 -5686 269749 -5652
rect 269737 -5692 269795 -5686
rect 269737 -5852 269795 -5846
rect 269737 -5886 269749 -5852
rect 269737 -5892 269795 -5886
rect 269924 -5901 269994 -5514
rect 270276 -5514 270310 -5513
rect 270698 -5513 270733 -5496
rect 271013 -5513 271048 -5496
rect 270698 -5514 270732 -5513
rect 270276 -5550 270346 -5514
rect 270106 -5581 270164 -5575
rect 270106 -5615 270118 -5581
rect 270293 -5584 270364 -5550
rect 270106 -5621 270164 -5615
rect 269924 -5935 269995 -5901
rect 270293 -5935 270363 -5584
rect 270475 -5652 270533 -5646
rect 270475 -5686 270487 -5652
rect 270475 -5692 270533 -5686
rect 270475 -5852 270533 -5846
rect 270475 -5886 270487 -5852
rect 270475 -5892 270533 -5886
rect 270662 -5901 270732 -5514
rect 271014 -5514 271048 -5513
rect 271436 -5513 271471 -5496
rect 271751 -5513 271786 -5496
rect 271436 -5514 271470 -5513
rect 271014 -5550 271084 -5514
rect 270844 -5581 270902 -5575
rect 270844 -5615 270856 -5581
rect 271031 -5584 271102 -5550
rect 270844 -5621 270902 -5615
rect 270662 -5935 270733 -5901
rect 271031 -5935 271101 -5584
rect 271213 -5652 271271 -5646
rect 271213 -5686 271225 -5652
rect 271213 -5692 271271 -5686
rect 271213 -5852 271271 -5846
rect 271213 -5886 271225 -5852
rect 271213 -5892 271271 -5886
rect 271400 -5901 271470 -5514
rect 271752 -5514 271786 -5513
rect 272174 -5513 272209 -5496
rect 272489 -5513 272524 -5496
rect 272174 -5514 272208 -5513
rect 271752 -5550 271822 -5514
rect 271582 -5581 271640 -5575
rect 271582 -5615 271594 -5581
rect 271769 -5584 271840 -5550
rect 271582 -5621 271640 -5615
rect 271400 -5935 271471 -5901
rect 271769 -5935 271839 -5584
rect 271951 -5652 272009 -5646
rect 271951 -5686 271963 -5652
rect 271951 -5692 272009 -5686
rect 271951 -5852 272009 -5846
rect 271951 -5886 271963 -5852
rect 271951 -5892 272009 -5886
rect 272138 -5901 272208 -5514
rect 272490 -5514 272524 -5513
rect 272912 -5513 272947 -5496
rect 273227 -5513 273262 -5496
rect 272912 -5514 272946 -5513
rect 272490 -5550 272560 -5514
rect 272320 -5581 272378 -5575
rect 272320 -5615 272332 -5581
rect 272507 -5584 272578 -5550
rect 272320 -5621 272378 -5615
rect 272138 -5935 272209 -5901
rect 272507 -5935 272577 -5584
rect 272689 -5652 272747 -5646
rect 272689 -5686 272701 -5652
rect 272689 -5692 272747 -5686
rect 272689 -5852 272747 -5846
rect 272689 -5886 272701 -5852
rect 272689 -5892 272747 -5886
rect 272876 -5901 272946 -5514
rect 273228 -5514 273262 -5513
rect 273650 -5513 273685 -5496
rect 273965 -5513 274000 -5496
rect 273650 -5514 273684 -5513
rect 273228 -5550 273298 -5514
rect 273058 -5581 273116 -5575
rect 273058 -5615 273070 -5581
rect 273245 -5584 273316 -5550
rect 273058 -5621 273116 -5615
rect 272876 -5935 272947 -5901
rect 273245 -5935 273315 -5584
rect 273427 -5652 273485 -5646
rect 273427 -5686 273439 -5652
rect 273427 -5692 273485 -5686
rect 273427 -5852 273485 -5846
rect 273427 -5886 273439 -5852
rect 273427 -5892 273485 -5886
rect 273614 -5901 273684 -5514
rect 273966 -5514 274000 -5513
rect 274388 -5513 274423 -5496
rect 274703 -5513 274738 -5496
rect 274388 -5514 274422 -5513
rect 273966 -5550 274036 -5514
rect 273796 -5581 273854 -5575
rect 273796 -5615 273808 -5581
rect 273983 -5584 274054 -5550
rect 273796 -5621 273854 -5615
rect 273614 -5935 273685 -5901
rect 273983 -5935 274053 -5584
rect 274165 -5652 274223 -5646
rect 274165 -5686 274177 -5652
rect 274165 -5692 274223 -5686
rect 274165 -5852 274223 -5846
rect 274165 -5886 274177 -5852
rect 274165 -5892 274223 -5886
rect 274352 -5901 274422 -5514
rect 274704 -5514 274738 -5513
rect 275126 -5513 275161 -5496
rect 275441 -5513 275476 -5496
rect 275126 -5514 275160 -5513
rect 274704 -5550 274774 -5514
rect 274534 -5581 274592 -5575
rect 274534 -5615 274546 -5581
rect 274721 -5584 274792 -5550
rect 274534 -5621 274592 -5615
rect 274352 -5935 274423 -5901
rect 274721 -5935 274791 -5584
rect 274903 -5652 274961 -5646
rect 274903 -5686 274915 -5652
rect 274903 -5692 274961 -5686
rect 274903 -5852 274961 -5846
rect 274903 -5886 274915 -5852
rect 274903 -5892 274961 -5886
rect 275090 -5901 275160 -5514
rect 275442 -5514 275476 -5513
rect 275864 -5513 275899 -5496
rect 276179 -5513 276214 -5496
rect 275864 -5514 275898 -5513
rect 275442 -5550 275512 -5514
rect 275272 -5581 275330 -5575
rect 275272 -5615 275284 -5581
rect 275459 -5584 275530 -5550
rect 275272 -5621 275330 -5615
rect 275090 -5935 275161 -5901
rect 275459 -5935 275529 -5584
rect 275641 -5652 275699 -5646
rect 275641 -5686 275653 -5652
rect 275641 -5692 275699 -5686
rect 275641 -5852 275699 -5846
rect 275641 -5886 275653 -5852
rect 275641 -5892 275699 -5886
rect 275828 -5901 275898 -5514
rect 276180 -5514 276214 -5513
rect 276602 -5513 276637 -5496
rect 276917 -5513 276952 -5496
rect 276602 -5514 276636 -5513
rect 276180 -5550 276250 -5514
rect 276010 -5581 276068 -5575
rect 276010 -5615 276022 -5581
rect 276197 -5584 276268 -5550
rect 276010 -5621 276068 -5615
rect 275828 -5935 275899 -5901
rect 276197 -5935 276267 -5584
rect 276379 -5652 276437 -5646
rect 276379 -5686 276391 -5652
rect 276379 -5692 276437 -5686
rect 276379 -5852 276437 -5846
rect 276379 -5886 276391 -5852
rect 276379 -5892 276437 -5886
rect 276566 -5901 276636 -5514
rect 276918 -5514 276952 -5513
rect 277340 -5513 277375 -5496
rect 277655 -5513 277690 -5496
rect 277340 -5514 277374 -5513
rect 276918 -5550 276988 -5514
rect 276748 -5581 276806 -5575
rect 276748 -5615 276760 -5581
rect 276935 -5584 277006 -5550
rect 276748 -5621 276806 -5615
rect 276566 -5935 276637 -5901
rect 276935 -5935 277005 -5584
rect 277117 -5652 277175 -5646
rect 277117 -5686 277129 -5652
rect 277117 -5692 277175 -5686
rect 277117 -5852 277175 -5846
rect 277117 -5886 277129 -5852
rect 277117 -5892 277175 -5886
rect 277304 -5901 277374 -5514
rect 277656 -5514 277690 -5513
rect 278078 -5513 278113 -5496
rect 278393 -5513 278428 -5496
rect 278078 -5514 278112 -5513
rect 277656 -5550 277726 -5514
rect 277486 -5581 277544 -5575
rect 277486 -5615 277498 -5581
rect 277673 -5584 277744 -5550
rect 277486 -5621 277544 -5615
rect 277304 -5935 277375 -5901
rect 277673 -5935 277743 -5584
rect 277855 -5652 277913 -5646
rect 277855 -5686 277867 -5652
rect 277855 -5692 277913 -5686
rect 277855 -5852 277913 -5846
rect 277855 -5886 277867 -5852
rect 277855 -5892 277913 -5886
rect 278042 -5901 278112 -5514
rect 278394 -5514 278428 -5513
rect 278816 -5513 278851 -5496
rect 279131 -5513 279166 -5496
rect 278816 -5514 278850 -5513
rect 278394 -5550 278464 -5514
rect 278224 -5581 278282 -5575
rect 278224 -5615 278236 -5581
rect 278411 -5584 278482 -5550
rect 278224 -5621 278282 -5615
rect 278042 -5935 278113 -5901
rect 278411 -5935 278481 -5584
rect 278593 -5652 278651 -5646
rect 278593 -5686 278605 -5652
rect 278593 -5692 278651 -5686
rect 278593 -5852 278651 -5846
rect 278593 -5886 278605 -5852
rect 278593 -5892 278651 -5886
rect 278780 -5901 278850 -5514
rect 279132 -5514 279166 -5513
rect 279554 -5513 279589 -5496
rect 279869 -5513 279904 -5496
rect 279554 -5514 279588 -5513
rect 279132 -5550 279202 -5514
rect 278962 -5581 279020 -5575
rect 278962 -5615 278974 -5581
rect 279149 -5584 279220 -5550
rect 278962 -5621 279020 -5615
rect 278780 -5935 278851 -5901
rect 279149 -5935 279219 -5584
rect 279331 -5652 279389 -5646
rect 279331 -5686 279343 -5652
rect 279331 -5692 279389 -5686
rect 279331 -5852 279389 -5846
rect 279331 -5886 279343 -5852
rect 279331 -5892 279389 -5886
rect 279518 -5901 279588 -5514
rect 279870 -5514 279904 -5513
rect 280292 -5513 280327 -5496
rect 280607 -5513 280642 -5496
rect 280292 -5514 280326 -5513
rect 279870 -5550 279940 -5514
rect 279700 -5581 279758 -5575
rect 279700 -5615 279712 -5581
rect 279887 -5584 279958 -5550
rect 279700 -5621 279758 -5615
rect 279518 -5935 279589 -5901
rect 279887 -5935 279957 -5584
rect 280069 -5652 280127 -5646
rect 280069 -5686 280081 -5652
rect 280069 -5692 280127 -5686
rect 280069 -5852 280127 -5846
rect 280069 -5886 280081 -5852
rect 280069 -5892 280127 -5886
rect 280256 -5901 280326 -5514
rect 280608 -5514 280642 -5513
rect 281030 -5513 281065 -5496
rect 281345 -5513 281380 -5496
rect 281030 -5514 281064 -5513
rect 280608 -5550 280678 -5514
rect 280438 -5581 280496 -5575
rect 280438 -5615 280450 -5581
rect 280625 -5584 280696 -5550
rect 280438 -5621 280496 -5615
rect 280256 -5935 280327 -5901
rect 280625 -5935 280695 -5584
rect 280807 -5652 280865 -5646
rect 280807 -5686 280819 -5652
rect 280807 -5692 280865 -5686
rect 280807 -5852 280865 -5846
rect 280807 -5886 280819 -5852
rect 280807 -5892 280865 -5886
rect 280994 -5901 281064 -5514
rect 281346 -5514 281380 -5513
rect 281768 -5513 281803 -5496
rect 282083 -5513 282118 -5496
rect 281768 -5514 281802 -5513
rect 281346 -5550 281416 -5514
rect 281176 -5581 281234 -5575
rect 281176 -5615 281188 -5581
rect 281363 -5584 281434 -5550
rect 281176 -5621 281234 -5615
rect 280994 -5935 281065 -5901
rect 281363 -5935 281433 -5584
rect 281545 -5652 281603 -5646
rect 281545 -5686 281557 -5652
rect 281545 -5692 281603 -5686
rect 281545 -5852 281603 -5846
rect 281545 -5886 281557 -5852
rect 281545 -5892 281603 -5886
rect 281732 -5901 281802 -5514
rect 282084 -5514 282118 -5513
rect 282506 -5513 282541 -5496
rect 282821 -5513 282856 -5496
rect 282506 -5514 282540 -5513
rect 282084 -5550 282154 -5514
rect 281914 -5581 281972 -5575
rect 281914 -5615 281926 -5581
rect 282101 -5584 282172 -5550
rect 281914 -5621 281972 -5615
rect 281732 -5935 281803 -5901
rect 282101 -5935 282171 -5584
rect 282283 -5652 282341 -5646
rect 282283 -5686 282295 -5652
rect 282283 -5692 282341 -5686
rect 282283 -5852 282341 -5846
rect 282283 -5886 282295 -5852
rect 282283 -5892 282341 -5886
rect 282470 -5901 282540 -5514
rect 282822 -5514 282856 -5513
rect 283244 -5513 283279 -5496
rect 283559 -5513 283594 -5496
rect 283244 -5514 283278 -5513
rect 282822 -5550 282892 -5514
rect 282652 -5581 282710 -5575
rect 282652 -5615 282664 -5581
rect 282839 -5584 282910 -5550
rect 282652 -5621 282710 -5615
rect 282470 -5935 282541 -5901
rect 282839 -5935 282909 -5584
rect 283021 -5652 283079 -5646
rect 283021 -5686 283033 -5652
rect 283021 -5692 283079 -5686
rect 283021 -5852 283079 -5846
rect 283021 -5886 283033 -5852
rect 283021 -5892 283079 -5886
rect 283208 -5901 283278 -5514
rect 283560 -5514 283594 -5513
rect 283982 -5513 284017 -5496
rect 284297 -5513 284332 -5496
rect 283982 -5514 284016 -5513
rect 283560 -5550 283630 -5514
rect 283390 -5581 283448 -5575
rect 283390 -5615 283402 -5581
rect 283577 -5584 283648 -5550
rect 283390 -5621 283448 -5615
rect 283208 -5935 283279 -5901
rect 283577 -5935 283647 -5584
rect 283759 -5652 283817 -5646
rect 283759 -5686 283771 -5652
rect 283759 -5692 283817 -5686
rect 283759 -5852 283817 -5846
rect 283759 -5886 283771 -5852
rect 283759 -5892 283817 -5886
rect 283946 -5901 284016 -5514
rect 284298 -5514 284332 -5513
rect 284720 -5513 284755 -5496
rect 285035 -5513 285070 -5496
rect 284720 -5514 284754 -5513
rect 284298 -5550 284368 -5514
rect 284128 -5581 284186 -5575
rect 284128 -5615 284140 -5581
rect 284315 -5584 284386 -5550
rect 284128 -5621 284186 -5615
rect 283946 -5935 284017 -5901
rect 284315 -5935 284385 -5584
rect 284497 -5652 284555 -5646
rect 284497 -5686 284509 -5652
rect 284497 -5692 284555 -5686
rect 284497 -5852 284555 -5846
rect 284497 -5886 284509 -5852
rect 284497 -5892 284555 -5886
rect 284684 -5901 284754 -5514
rect 285036 -5514 285070 -5513
rect 285458 -5513 285493 -5496
rect 285773 -5513 285808 -5496
rect 285458 -5514 285492 -5513
rect 285036 -5550 285106 -5514
rect 284866 -5581 284924 -5575
rect 284866 -5615 284878 -5581
rect 285053 -5584 285124 -5550
rect 284866 -5621 284924 -5615
rect 284684 -5935 284755 -5901
rect 285053 -5935 285123 -5584
rect 285235 -5652 285293 -5646
rect 285235 -5686 285247 -5652
rect 285235 -5692 285293 -5686
rect 285235 -5852 285293 -5846
rect 285235 -5886 285247 -5852
rect 285235 -5892 285293 -5886
rect 285422 -5901 285492 -5514
rect 285774 -5514 285808 -5513
rect 286196 -5513 286231 -5496
rect 286511 -5513 286546 -5496
rect 286196 -5514 286230 -5513
rect 285774 -5550 285844 -5514
rect 285604 -5581 285662 -5575
rect 285604 -5615 285616 -5581
rect 285791 -5584 285862 -5550
rect 285604 -5621 285662 -5615
rect 285422 -5935 285493 -5901
rect 285791 -5935 285861 -5584
rect 285973 -5652 286031 -5646
rect 285973 -5686 285985 -5652
rect 285973 -5692 286031 -5686
rect 285973 -5852 286031 -5846
rect 285973 -5886 285985 -5852
rect 285973 -5892 286031 -5886
rect 286160 -5901 286230 -5514
rect 286512 -5514 286546 -5513
rect 286934 -5513 286969 -5496
rect 287249 -5513 287284 -5496
rect 286934 -5514 286968 -5513
rect 286512 -5550 286582 -5514
rect 286342 -5581 286400 -5575
rect 286342 -5615 286354 -5581
rect 286529 -5584 286600 -5550
rect 286342 -5621 286400 -5615
rect 286160 -5935 286231 -5901
rect 286529 -5935 286599 -5584
rect 286711 -5652 286769 -5646
rect 286711 -5686 286723 -5652
rect 286711 -5692 286769 -5686
rect 286711 -5852 286769 -5846
rect 286711 -5886 286723 -5852
rect 286711 -5892 286769 -5886
rect 286898 -5901 286968 -5514
rect 287250 -5514 287284 -5513
rect 287672 -5513 287707 -5496
rect 287987 -5513 288022 -5496
rect 287672 -5514 287706 -5513
rect 287250 -5550 287320 -5514
rect 287080 -5581 287138 -5575
rect 287080 -5615 287092 -5581
rect 287267 -5584 287338 -5550
rect 287080 -5621 287138 -5615
rect 286898 -5935 286969 -5901
rect 287267 -5935 287337 -5584
rect 287449 -5652 287507 -5646
rect 287449 -5686 287461 -5652
rect 287449 -5692 287507 -5686
rect 287449 -5852 287507 -5846
rect 287449 -5886 287461 -5852
rect 287449 -5892 287507 -5886
rect 287636 -5901 287706 -5514
rect 287988 -5514 288022 -5513
rect 288410 -5513 288445 -5496
rect 288725 -5513 288760 -5496
rect 288410 -5514 288444 -5513
rect 287988 -5550 288058 -5514
rect 287818 -5581 287876 -5575
rect 287818 -5615 287830 -5581
rect 288005 -5584 288076 -5550
rect 287818 -5621 287876 -5615
rect 287636 -5935 287707 -5901
rect 288005 -5935 288075 -5584
rect 288187 -5652 288245 -5646
rect 288187 -5686 288199 -5652
rect 288187 -5692 288245 -5686
rect 288187 -5852 288245 -5846
rect 288187 -5886 288199 -5852
rect 288187 -5892 288245 -5886
rect 288374 -5901 288444 -5514
rect 288726 -5514 288760 -5513
rect 289148 -5513 289183 -5496
rect 289463 -5513 289498 -5496
rect 289148 -5514 289182 -5513
rect 288726 -5550 288796 -5514
rect 288556 -5581 288614 -5575
rect 288556 -5615 288568 -5581
rect 288743 -5584 288814 -5550
rect 288556 -5621 288614 -5615
rect 288374 -5935 288445 -5901
rect 288743 -5935 288813 -5584
rect 288925 -5652 288983 -5646
rect 288925 -5686 288937 -5652
rect 288925 -5692 288983 -5686
rect 288925 -5852 288983 -5846
rect 288925 -5886 288937 -5852
rect 288925 -5892 288983 -5886
rect 289112 -5901 289182 -5514
rect 289464 -5514 289498 -5513
rect 289886 -5513 289921 -5496
rect 290201 -5513 290236 -5496
rect 289886 -5514 289920 -5513
rect 289464 -5550 289534 -5514
rect 289294 -5581 289352 -5575
rect 289294 -5615 289306 -5581
rect 289481 -5584 289552 -5550
rect 289294 -5621 289352 -5615
rect 289112 -5935 289183 -5901
rect 289481 -5935 289551 -5584
rect 289663 -5652 289721 -5646
rect 289663 -5686 289675 -5652
rect 289663 -5692 289721 -5686
rect 289663 -5852 289721 -5846
rect 289663 -5886 289675 -5852
rect 289663 -5892 289721 -5886
rect 289850 -5901 289920 -5514
rect 290202 -5514 290236 -5513
rect 290624 -5513 290659 -5496
rect 290939 -5513 290974 -5496
rect 290624 -5514 290658 -5513
rect 290202 -5550 290272 -5514
rect 290032 -5581 290090 -5575
rect 290032 -5615 290044 -5581
rect 290219 -5584 290290 -5550
rect 290032 -5621 290090 -5615
rect 289850 -5935 289921 -5901
rect 290219 -5935 290289 -5584
rect 290401 -5652 290459 -5646
rect 290401 -5686 290413 -5652
rect 290401 -5692 290459 -5686
rect 290401 -5852 290459 -5846
rect 290401 -5886 290413 -5852
rect 290401 -5892 290459 -5886
rect 290588 -5901 290658 -5514
rect 290940 -5514 290974 -5513
rect 291362 -5513 291397 -5496
rect 291677 -5513 291712 -5496
rect 291362 -5514 291396 -5513
rect 290940 -5550 291010 -5514
rect 290770 -5581 290828 -5575
rect 290770 -5615 290782 -5581
rect 290957 -5584 291028 -5550
rect 290770 -5621 290828 -5615
rect 290588 -5935 290659 -5901
rect 290957 -5935 291027 -5584
rect 291139 -5652 291197 -5646
rect 291139 -5686 291151 -5652
rect 291139 -5692 291197 -5686
rect 291139 -5852 291197 -5846
rect 291139 -5886 291151 -5852
rect 291139 -5892 291197 -5886
rect 291326 -5901 291396 -5514
rect 291678 -5514 291712 -5513
rect 292100 -5513 292135 -5496
rect 292415 -5513 292450 -5496
rect 292100 -5514 292134 -5513
rect 291678 -5550 291748 -5514
rect 291508 -5581 291566 -5575
rect 291508 -5615 291520 -5581
rect 291695 -5584 291766 -5550
rect 291508 -5621 291566 -5615
rect 291326 -5935 291397 -5901
rect 291695 -5935 291765 -5584
rect 291877 -5652 291935 -5646
rect 291877 -5686 291889 -5652
rect 291877 -5692 291935 -5686
rect 291877 -5852 291935 -5846
rect 291877 -5886 291889 -5852
rect 291877 -5892 291935 -5886
rect 292064 -5901 292134 -5514
rect 292416 -5514 292450 -5513
rect 292838 -5513 292873 -5496
rect 293153 -5513 293188 -5496
rect 292838 -5514 292872 -5513
rect 292416 -5550 292486 -5514
rect 292246 -5581 292304 -5575
rect 292246 -5615 292258 -5581
rect 292433 -5584 292504 -5550
rect 292246 -5621 292304 -5615
rect 292064 -5935 292135 -5901
rect 292433 -5935 292503 -5584
rect 292615 -5652 292673 -5646
rect 292615 -5686 292627 -5652
rect 292615 -5692 292673 -5686
rect 292615 -5852 292673 -5846
rect 292615 -5886 292627 -5852
rect 292615 -5892 292673 -5886
rect 292802 -5901 292872 -5514
rect 293154 -5514 293188 -5513
rect 293576 -5513 293611 -5496
rect 293891 -5513 293926 -5496
rect 293576 -5514 293610 -5513
rect 293154 -5550 293224 -5514
rect 292984 -5581 293042 -5575
rect 292984 -5615 292996 -5581
rect 293171 -5584 293242 -5550
rect 292984 -5621 293042 -5615
rect 292802 -5935 292873 -5901
rect 293171 -5935 293241 -5584
rect 293353 -5652 293411 -5646
rect 293353 -5686 293365 -5652
rect 293353 -5692 293411 -5686
rect 293353 -5852 293411 -5846
rect 293353 -5886 293365 -5852
rect 293353 -5892 293411 -5886
rect 293540 -5901 293610 -5514
rect 293892 -5514 293926 -5513
rect 294314 -5513 294349 -5496
rect 294629 -5513 294664 -5496
rect 294314 -5514 294348 -5513
rect 293892 -5550 293962 -5514
rect 293722 -5581 293780 -5575
rect 293722 -5615 293734 -5581
rect 293909 -5584 293980 -5550
rect 293722 -5621 293780 -5615
rect 293540 -5935 293611 -5901
rect 293909 -5935 293979 -5584
rect 294091 -5652 294149 -5646
rect 294091 -5686 294103 -5652
rect 294091 -5692 294149 -5686
rect 294091 -5852 294149 -5846
rect 294091 -5886 294103 -5852
rect 294091 -5892 294149 -5886
rect 294278 -5901 294348 -5514
rect 294630 -5514 294664 -5513
rect 295052 -5513 295087 -5496
rect 295367 -5513 295402 -5496
rect 295052 -5514 295086 -5513
rect 294630 -5550 294700 -5514
rect 294460 -5581 294518 -5575
rect 294460 -5615 294472 -5581
rect 294647 -5584 294718 -5550
rect 294460 -5621 294518 -5615
rect 294278 -5935 294349 -5901
rect 294647 -5935 294717 -5584
rect 294829 -5652 294887 -5646
rect 294829 -5686 294841 -5652
rect 294829 -5692 294887 -5686
rect 294829 -5852 294887 -5846
rect 294829 -5886 294841 -5852
rect 294829 -5892 294887 -5886
rect 295016 -5901 295086 -5514
rect 295368 -5514 295402 -5513
rect 295790 -5513 295825 -5496
rect 296105 -5513 296140 -5496
rect 295790 -5514 295824 -5513
rect 295368 -5550 295438 -5514
rect 295198 -5581 295256 -5575
rect 295198 -5615 295210 -5581
rect 295385 -5584 295456 -5550
rect 295198 -5621 295256 -5615
rect 295016 -5935 295087 -5901
rect 295385 -5935 295455 -5584
rect 295567 -5652 295625 -5646
rect 295567 -5686 295579 -5652
rect 295567 -5692 295625 -5686
rect 295567 -5852 295625 -5846
rect 295567 -5886 295579 -5852
rect 295567 -5892 295625 -5886
rect 295754 -5901 295824 -5514
rect 296106 -5514 296140 -5513
rect 296528 -5513 296563 -5496
rect 296843 -5513 296878 -5496
rect 296528 -5514 296562 -5513
rect 296106 -5550 296176 -5514
rect 295936 -5581 295994 -5575
rect 295936 -5615 295948 -5581
rect 296123 -5584 296194 -5550
rect 295936 -5621 295994 -5615
rect 295754 -5935 295825 -5901
rect 296123 -5935 296193 -5584
rect 296305 -5652 296363 -5646
rect 296305 -5686 296317 -5652
rect 296305 -5692 296363 -5686
rect 296305 -5852 296363 -5846
rect 296305 -5886 296317 -5852
rect 296305 -5892 296363 -5886
rect 296492 -5901 296562 -5514
rect 296844 -5514 296878 -5513
rect 297266 -5513 297301 -5496
rect 297581 -5513 297616 -5496
rect 297266 -5514 297300 -5513
rect 296844 -5550 296914 -5514
rect 296674 -5581 296732 -5575
rect 296674 -5615 296686 -5581
rect 296861 -5584 296932 -5550
rect 296674 -5621 296732 -5615
rect 296492 -5935 296563 -5901
rect 296861 -5935 296931 -5584
rect 297043 -5652 297101 -5646
rect 297043 -5686 297055 -5652
rect 297043 -5692 297101 -5686
rect 297043 -5852 297101 -5846
rect 297043 -5886 297055 -5852
rect 297043 -5892 297101 -5886
rect 297230 -5901 297300 -5514
rect 297582 -5514 297616 -5513
rect 298004 -5513 298039 -5496
rect 298319 -5513 298354 -5496
rect 298004 -5514 298038 -5513
rect 297582 -5550 297652 -5514
rect 297412 -5581 297470 -5575
rect 297412 -5615 297424 -5581
rect 297599 -5584 297670 -5550
rect 297412 -5621 297470 -5615
rect 297230 -5935 297301 -5901
rect 297599 -5935 297669 -5584
rect 297781 -5652 297839 -5646
rect 297781 -5686 297793 -5652
rect 297781 -5692 297839 -5686
rect 297781 -5852 297839 -5846
rect 297781 -5886 297793 -5852
rect 297781 -5892 297839 -5886
rect 297968 -5901 298038 -5514
rect 298320 -5514 298354 -5513
rect 298742 -5513 298777 -5496
rect 299057 -5513 299092 -5496
rect 298742 -5514 298776 -5513
rect 298320 -5550 298390 -5514
rect 298150 -5581 298208 -5575
rect 298150 -5615 298162 -5581
rect 298337 -5584 298408 -5550
rect 298150 -5621 298208 -5615
rect 297968 -5935 298039 -5901
rect 298337 -5935 298407 -5584
rect 298519 -5652 298577 -5646
rect 298519 -5686 298531 -5652
rect 298519 -5692 298577 -5686
rect 298519 -5852 298577 -5846
rect 298519 -5886 298531 -5852
rect 298519 -5892 298577 -5886
rect 298706 -5901 298776 -5514
rect 299058 -5514 299092 -5513
rect 299480 -5513 299515 -5496
rect 299795 -5513 299830 -5496
rect 299480 -5514 299514 -5513
rect 299058 -5550 299128 -5514
rect 298888 -5581 298946 -5575
rect 298888 -5615 298900 -5581
rect 299075 -5584 299146 -5550
rect 298888 -5621 298946 -5615
rect 298706 -5935 298777 -5901
rect 299075 -5935 299145 -5584
rect 299257 -5652 299315 -5646
rect 299257 -5686 299269 -5652
rect 299257 -5692 299315 -5686
rect 299257 -5852 299315 -5846
rect 299257 -5886 299269 -5852
rect 299257 -5892 299315 -5886
rect 299444 -5901 299514 -5514
rect 299796 -5514 299830 -5513
rect 300218 -5513 300253 -5496
rect 300533 -5513 300568 -5496
rect 300218 -5514 300252 -5513
rect 299796 -5550 299866 -5514
rect 299626 -5581 299684 -5575
rect 299626 -5615 299638 -5581
rect 299813 -5584 299884 -5550
rect 299626 -5621 299684 -5615
rect 299444 -5935 299515 -5901
rect 299813 -5935 299883 -5584
rect 299995 -5652 300053 -5646
rect 299995 -5686 300007 -5652
rect 299995 -5692 300053 -5686
rect 299995 -5852 300053 -5846
rect 299995 -5886 300007 -5852
rect 299995 -5892 300053 -5886
rect 300182 -5901 300252 -5514
rect 300534 -5514 300568 -5513
rect 300956 -5513 300991 -5496
rect 301271 -5513 301306 -5496
rect 300956 -5514 300990 -5513
rect 300534 -5550 300604 -5514
rect 300364 -5581 300422 -5575
rect 300364 -5615 300376 -5581
rect 300551 -5584 300622 -5550
rect 300364 -5621 300422 -5615
rect 300182 -5935 300253 -5901
rect 300551 -5935 300621 -5584
rect 300733 -5652 300791 -5646
rect 300733 -5686 300745 -5652
rect 300733 -5692 300791 -5686
rect 300733 -5852 300791 -5846
rect 300733 -5886 300745 -5852
rect 300733 -5892 300791 -5886
rect 300920 -5901 300990 -5514
rect 301272 -5514 301306 -5513
rect 301694 -5513 301729 -5496
rect 302009 -5513 302044 -5496
rect 301694 -5514 301728 -5513
rect 301272 -5550 301342 -5514
rect 301102 -5581 301160 -5575
rect 301102 -5615 301114 -5581
rect 301289 -5584 301360 -5550
rect 301102 -5621 301160 -5615
rect 300920 -5935 300991 -5901
rect 301289 -5935 301359 -5584
rect 301471 -5652 301529 -5646
rect 301471 -5686 301483 -5652
rect 301471 -5692 301529 -5686
rect 301471 -5852 301529 -5846
rect 301471 -5886 301483 -5852
rect 301471 -5892 301529 -5886
rect 301658 -5901 301728 -5514
rect 302010 -5514 302044 -5513
rect 302432 -5513 302467 -5496
rect 302747 -5513 302782 -5496
rect 302432 -5514 302466 -5513
rect 302010 -5550 302080 -5514
rect 301840 -5581 301898 -5575
rect 301840 -5615 301852 -5581
rect 302027 -5584 302098 -5550
rect 301840 -5621 301898 -5615
rect 301658 -5935 301729 -5901
rect 302027 -5935 302097 -5584
rect 302209 -5652 302267 -5646
rect 302209 -5686 302221 -5652
rect 302209 -5692 302267 -5686
rect 302209 -5852 302267 -5846
rect 302209 -5886 302221 -5852
rect 302209 -5892 302267 -5886
rect 302396 -5901 302466 -5514
rect 302748 -5514 302782 -5513
rect 303170 -5513 303205 -5496
rect 303485 -5513 303520 -5496
rect 303170 -5514 303204 -5513
rect 302748 -5550 302818 -5514
rect 302578 -5581 302636 -5575
rect 302578 -5615 302590 -5581
rect 302765 -5584 302836 -5550
rect 302578 -5621 302636 -5615
rect 302396 -5935 302467 -5901
rect 302765 -5935 302835 -5584
rect 302947 -5652 303005 -5646
rect 302947 -5686 302959 -5652
rect 302947 -5692 303005 -5686
rect 302947 -5852 303005 -5846
rect 302947 -5886 302959 -5852
rect 302947 -5892 303005 -5886
rect 303134 -5901 303204 -5514
rect 303486 -5514 303520 -5513
rect 303908 -5513 303943 -5496
rect 304223 -5513 304258 -5496
rect 303908 -5514 303942 -5513
rect 303486 -5550 303556 -5514
rect 303316 -5581 303374 -5575
rect 303316 -5615 303328 -5581
rect 303503 -5584 303574 -5550
rect 303316 -5621 303374 -5615
rect 303134 -5935 303205 -5901
rect 303503 -5935 303573 -5584
rect 303685 -5652 303743 -5646
rect 303685 -5686 303697 -5652
rect 303685 -5692 303743 -5686
rect 303685 -5852 303743 -5846
rect 303685 -5886 303697 -5852
rect 303685 -5892 303743 -5886
rect 303872 -5901 303942 -5514
rect 304224 -5514 304258 -5513
rect 304646 -5513 304681 -5496
rect 304961 -5513 304996 -5496
rect 304646 -5514 304680 -5513
rect 304224 -5550 304294 -5514
rect 304054 -5581 304112 -5575
rect 304054 -5615 304066 -5581
rect 304241 -5584 304312 -5550
rect 304054 -5621 304112 -5615
rect 303872 -5935 303943 -5901
rect 304241 -5935 304311 -5584
rect 304423 -5652 304481 -5646
rect 304423 -5686 304435 -5652
rect 304423 -5692 304481 -5686
rect 304423 -5852 304481 -5846
rect 304423 -5886 304435 -5852
rect 304423 -5892 304481 -5886
rect 304610 -5901 304680 -5514
rect 304962 -5514 304996 -5513
rect 305384 -5513 305419 -5496
rect 305699 -5513 305734 -5496
rect 305384 -5514 305418 -5513
rect 304962 -5550 305032 -5514
rect 304792 -5581 304850 -5575
rect 304792 -5615 304804 -5581
rect 304979 -5584 305050 -5550
rect 304792 -5621 304850 -5615
rect 304610 -5935 304681 -5901
rect 304979 -5935 305049 -5584
rect 305161 -5652 305219 -5646
rect 305161 -5686 305173 -5652
rect 305161 -5692 305219 -5686
rect 305161 -5852 305219 -5846
rect 305161 -5886 305173 -5852
rect 305161 -5892 305219 -5886
rect 305348 -5901 305418 -5514
rect 305700 -5514 305734 -5513
rect 306122 -5513 306157 -5496
rect 306437 -5513 306472 -5496
rect 306122 -5514 306156 -5513
rect 305700 -5550 305770 -5514
rect 305530 -5581 305588 -5575
rect 305530 -5615 305542 -5581
rect 305717 -5584 305788 -5550
rect 305530 -5621 305588 -5615
rect 305348 -5935 305419 -5901
rect 305717 -5935 305787 -5584
rect 305899 -5652 305957 -5646
rect 305899 -5686 305911 -5652
rect 305899 -5692 305957 -5686
rect 305899 -5852 305957 -5846
rect 305899 -5886 305911 -5852
rect 305899 -5892 305957 -5886
rect 306086 -5901 306156 -5514
rect 306438 -5514 306472 -5513
rect 306860 -5513 306895 -5496
rect 307175 -5513 307210 -5496
rect 306860 -5514 306894 -5513
rect 306438 -5550 306508 -5514
rect 306268 -5581 306326 -5575
rect 306268 -5615 306280 -5581
rect 306455 -5584 306526 -5550
rect 306268 -5621 306326 -5615
rect 306086 -5935 306157 -5901
rect 306455 -5935 306525 -5584
rect 306637 -5652 306695 -5646
rect 306637 -5686 306649 -5652
rect 306637 -5692 306695 -5686
rect 306637 -5852 306695 -5846
rect 306637 -5886 306649 -5852
rect 306637 -5892 306695 -5886
rect 306824 -5901 306894 -5514
rect 307176 -5514 307210 -5513
rect 307598 -5513 307633 -5496
rect 307913 -5513 307948 -5496
rect 307598 -5514 307632 -5513
rect 307176 -5550 307246 -5514
rect 307006 -5581 307064 -5575
rect 307006 -5615 307018 -5581
rect 307193 -5584 307264 -5550
rect 307006 -5621 307064 -5615
rect 306824 -5935 306895 -5901
rect 307193 -5935 307263 -5584
rect 307375 -5652 307433 -5646
rect 307375 -5686 307387 -5652
rect 307375 -5692 307433 -5686
rect 307375 -5852 307433 -5846
rect 307375 -5886 307387 -5852
rect 307375 -5892 307433 -5886
rect 307562 -5901 307632 -5514
rect 307914 -5514 307948 -5513
rect 308336 -5513 308371 -5496
rect 308651 -5513 308686 -5496
rect 308336 -5514 308370 -5513
rect 307914 -5550 307984 -5514
rect 307744 -5581 307802 -5575
rect 307744 -5615 307756 -5581
rect 307931 -5584 308002 -5550
rect 307744 -5621 307802 -5615
rect 307562 -5935 307633 -5901
rect 307931 -5935 308001 -5584
rect 308113 -5652 308171 -5646
rect 308113 -5686 308125 -5652
rect 308113 -5692 308171 -5686
rect 308113 -5852 308171 -5846
rect 308113 -5886 308125 -5852
rect 308113 -5892 308171 -5886
rect 308300 -5901 308370 -5514
rect 308652 -5514 308686 -5513
rect 309074 -5513 309109 -5496
rect 309389 -5513 309424 -5496
rect 309074 -5514 309108 -5513
rect 308652 -5550 308722 -5514
rect 308482 -5581 308540 -5575
rect 308482 -5615 308494 -5581
rect 308669 -5584 308740 -5550
rect 308482 -5621 308540 -5615
rect 308300 -5935 308371 -5901
rect 308669 -5935 308739 -5584
rect 308851 -5652 308909 -5646
rect 308851 -5686 308863 -5652
rect 308851 -5692 308909 -5686
rect 308851 -5852 308909 -5846
rect 308851 -5886 308863 -5852
rect 308851 -5892 308909 -5886
rect 309038 -5901 309108 -5514
rect 309390 -5514 309424 -5513
rect 309812 -5513 309847 -5496
rect 310127 -5513 310162 -5496
rect 309812 -5514 309846 -5513
rect 309390 -5550 309460 -5514
rect 309220 -5581 309278 -5575
rect 309220 -5615 309232 -5581
rect 309407 -5584 309478 -5550
rect 309220 -5621 309278 -5615
rect 309038 -5935 309109 -5901
rect 309407 -5935 309477 -5584
rect 309589 -5652 309647 -5646
rect 309589 -5686 309601 -5652
rect 309589 -5692 309647 -5686
rect 309589 -5852 309647 -5846
rect 309589 -5886 309601 -5852
rect 309589 -5892 309647 -5886
rect 309776 -5901 309846 -5514
rect 310128 -5514 310162 -5513
rect 310550 -5513 310585 -5496
rect 310865 -5513 310900 -5496
rect 310550 -5514 310584 -5513
rect 310128 -5550 310198 -5514
rect 309958 -5581 310016 -5575
rect 309958 -5615 309970 -5581
rect 310145 -5584 310216 -5550
rect 309958 -5621 310016 -5615
rect 309776 -5935 309847 -5901
rect 310145 -5935 310215 -5584
rect 310327 -5652 310385 -5646
rect 310327 -5686 310339 -5652
rect 310327 -5692 310385 -5686
rect 310327 -5852 310385 -5846
rect 310327 -5886 310339 -5852
rect 310327 -5892 310385 -5886
rect 310514 -5901 310584 -5514
rect 310866 -5514 310900 -5513
rect 311288 -5513 311323 -5496
rect 311603 -5513 311638 -5496
rect 311288 -5514 311322 -5513
rect 310866 -5550 310936 -5514
rect 310696 -5581 310754 -5575
rect 310696 -5615 310708 -5581
rect 310883 -5584 310954 -5550
rect 310696 -5621 310754 -5615
rect 310514 -5935 310585 -5901
rect 310883 -5935 310953 -5584
rect 311065 -5652 311123 -5646
rect 311065 -5686 311077 -5652
rect 311065 -5692 311123 -5686
rect 311065 -5852 311123 -5846
rect 311065 -5886 311077 -5852
rect 311065 -5892 311123 -5886
rect 311252 -5901 311322 -5514
rect 311604 -5514 311638 -5513
rect 312026 -5513 312061 -5496
rect 312341 -5513 312376 -5496
rect 312026 -5514 312060 -5513
rect 311604 -5550 311674 -5514
rect 311434 -5581 311492 -5575
rect 311434 -5615 311446 -5581
rect 311621 -5584 311692 -5550
rect 311434 -5621 311492 -5615
rect 311252 -5935 311323 -5901
rect 311621 -5935 311691 -5584
rect 311803 -5652 311861 -5646
rect 311803 -5686 311815 -5652
rect 311803 -5692 311861 -5686
rect 311803 -5852 311861 -5846
rect 311803 -5886 311815 -5852
rect 311803 -5892 311861 -5886
rect 311990 -5901 312060 -5514
rect 312342 -5514 312376 -5513
rect 312764 -5513 312799 -5496
rect 313079 -5513 313114 -5496
rect 312764 -5514 312798 -5513
rect 312342 -5550 312412 -5514
rect 312172 -5581 312230 -5575
rect 312172 -5615 312184 -5581
rect 312359 -5584 312430 -5550
rect 312172 -5621 312230 -5615
rect 311990 -5935 312061 -5901
rect 312359 -5935 312429 -5584
rect 312541 -5652 312599 -5646
rect 312541 -5686 312553 -5652
rect 312541 -5692 312599 -5686
rect 312541 -5852 312599 -5846
rect 312541 -5886 312553 -5852
rect 312541 -5892 312599 -5886
rect 312728 -5901 312798 -5514
rect 313080 -5514 313114 -5513
rect 313502 -5513 313537 -5496
rect 313817 -5513 313852 -5496
rect 313502 -5514 313536 -5513
rect 313080 -5550 313150 -5514
rect 312910 -5581 312968 -5575
rect 312910 -5615 312922 -5581
rect 313097 -5584 313168 -5550
rect 312910 -5621 312968 -5615
rect 312728 -5935 312799 -5901
rect 313097 -5935 313167 -5584
rect 313279 -5652 313337 -5646
rect 313279 -5686 313291 -5652
rect 313279 -5692 313337 -5686
rect 313279 -5852 313337 -5846
rect 313279 -5886 313291 -5852
rect 313279 -5892 313337 -5886
rect 313466 -5901 313536 -5514
rect 313818 -5514 313852 -5513
rect 314240 -5513 314275 -5496
rect 314555 -5513 314590 -5496
rect 314240 -5514 314274 -5513
rect 313818 -5550 313888 -5514
rect 313648 -5581 313706 -5575
rect 313648 -5615 313660 -5581
rect 313835 -5584 313906 -5550
rect 313648 -5621 313706 -5615
rect 313466 -5935 313537 -5901
rect 313835 -5935 313905 -5584
rect 314017 -5652 314075 -5646
rect 314017 -5686 314029 -5652
rect 314017 -5692 314075 -5686
rect 314017 -5852 314075 -5846
rect 314017 -5886 314029 -5852
rect 314017 -5892 314075 -5886
rect 314204 -5901 314274 -5514
rect 314556 -5514 314590 -5513
rect 314978 -5513 315013 -5496
rect 315293 -5513 315328 -5496
rect 314978 -5514 315012 -5513
rect 314556 -5550 314626 -5514
rect 314386 -5581 314444 -5575
rect 314386 -5615 314398 -5581
rect 314573 -5584 314644 -5550
rect 314386 -5621 314444 -5615
rect 314204 -5935 314275 -5901
rect 314573 -5935 314643 -5584
rect 314755 -5652 314813 -5646
rect 314755 -5686 314767 -5652
rect 314755 -5692 314813 -5686
rect 314755 -5852 314813 -5846
rect 314755 -5886 314767 -5852
rect 314755 -5892 314813 -5886
rect 314942 -5901 315012 -5514
rect 315294 -5514 315328 -5513
rect 315716 -5513 315751 -5496
rect 316031 -5513 316066 -5496
rect 315716 -5514 315750 -5513
rect 315294 -5550 315364 -5514
rect 315124 -5581 315182 -5575
rect 315124 -5615 315136 -5581
rect 315311 -5584 315382 -5550
rect 315124 -5621 315182 -5615
rect 314942 -5935 315013 -5901
rect 315311 -5935 315381 -5584
rect 315493 -5652 315551 -5646
rect 315493 -5686 315505 -5652
rect 315493 -5692 315551 -5686
rect 315493 -5852 315551 -5846
rect 315493 -5886 315505 -5852
rect 315493 -5892 315551 -5886
rect 315680 -5901 315750 -5514
rect 316032 -5514 316066 -5513
rect 316454 -5513 316489 -5496
rect 316769 -5513 316804 -5496
rect 316454 -5514 316488 -5513
rect 316032 -5550 316102 -5514
rect 315862 -5581 315920 -5575
rect 315862 -5615 315874 -5581
rect 316049 -5584 316120 -5550
rect 315862 -5621 315920 -5615
rect 315680 -5935 315751 -5901
rect 316049 -5935 316119 -5584
rect 316231 -5652 316289 -5646
rect 316231 -5686 316243 -5652
rect 316231 -5692 316289 -5686
rect 316231 -5852 316289 -5846
rect 316231 -5886 316243 -5852
rect 316231 -5892 316289 -5886
rect 316418 -5901 316488 -5514
rect 316770 -5514 316804 -5513
rect 317192 -5513 317227 -5496
rect 317507 -5513 317542 -5496
rect 317192 -5514 317226 -5513
rect 316770 -5550 316840 -5514
rect 316600 -5581 316658 -5575
rect 316600 -5615 316612 -5581
rect 316787 -5584 316858 -5550
rect 316600 -5621 316658 -5615
rect 316418 -5935 316489 -5901
rect 316787 -5935 316857 -5584
rect 316969 -5652 317027 -5646
rect 316969 -5686 316981 -5652
rect 316969 -5692 317027 -5686
rect 316969 -5852 317027 -5846
rect 316969 -5886 316981 -5852
rect 316969 -5892 317027 -5886
rect 317156 -5901 317226 -5514
rect 317508 -5514 317542 -5513
rect 317930 -5513 317965 -5496
rect 318245 -5513 318280 -5496
rect 317930 -5514 317964 -5513
rect 317508 -5550 317578 -5514
rect 317338 -5581 317396 -5575
rect 317338 -5615 317350 -5581
rect 317525 -5584 317596 -5550
rect 317338 -5621 317396 -5615
rect 317156 -5935 317227 -5901
rect 317525 -5935 317595 -5584
rect 317707 -5652 317765 -5646
rect 317707 -5686 317719 -5652
rect 317707 -5692 317765 -5686
rect 317707 -5852 317765 -5846
rect 317707 -5886 317719 -5852
rect 317707 -5892 317765 -5886
rect 317894 -5901 317964 -5514
rect 318246 -5514 318280 -5513
rect 318668 -5513 318703 -5496
rect 318983 -5513 319018 -5496
rect 318668 -5514 318702 -5513
rect 318246 -5550 318316 -5514
rect 318076 -5581 318134 -5575
rect 318076 -5615 318088 -5581
rect 318263 -5584 318334 -5550
rect 318076 -5621 318134 -5615
rect 317894 -5935 317965 -5901
rect 318263 -5935 318333 -5584
rect 318445 -5652 318503 -5646
rect 318445 -5686 318457 -5652
rect 318445 -5692 318503 -5686
rect 318445 -5852 318503 -5846
rect 318445 -5886 318457 -5852
rect 318445 -5892 318503 -5886
rect 318632 -5901 318702 -5514
rect 318984 -5514 319018 -5513
rect 319406 -5513 319441 -5496
rect 319721 -5513 319756 -5496
rect 319406 -5514 319440 -5513
rect 318984 -5550 319054 -5514
rect 318814 -5581 318872 -5575
rect 318814 -5615 318826 -5581
rect 319001 -5584 319072 -5550
rect 318814 -5621 318872 -5615
rect 318632 -5935 318703 -5901
rect 319001 -5935 319071 -5584
rect 319183 -5652 319241 -5646
rect 319183 -5686 319195 -5652
rect 319183 -5692 319241 -5686
rect 319183 -5852 319241 -5846
rect 319183 -5886 319195 -5852
rect 319183 -5892 319241 -5886
rect 319370 -5901 319440 -5514
rect 319722 -5514 319756 -5513
rect 320144 -5513 320179 -5496
rect 320459 -5513 320494 -5496
rect 320144 -5514 320178 -5513
rect 319722 -5550 319792 -5514
rect 319552 -5581 319610 -5575
rect 319552 -5615 319564 -5581
rect 319739 -5584 319810 -5550
rect 319552 -5621 319610 -5615
rect 319370 -5935 319441 -5901
rect 319739 -5935 319809 -5584
rect 319921 -5652 319979 -5646
rect 319921 -5686 319933 -5652
rect 319921 -5692 319979 -5686
rect 319921 -5852 319979 -5846
rect 319921 -5886 319933 -5852
rect 319921 -5892 319979 -5886
rect 320108 -5901 320178 -5514
rect 320460 -5514 320494 -5513
rect 320882 -5513 320917 -5496
rect 321197 -5513 321232 -5496
rect 320882 -5514 320916 -5513
rect 320460 -5550 320530 -5514
rect 320290 -5581 320348 -5575
rect 320290 -5615 320302 -5581
rect 320477 -5584 320548 -5550
rect 320290 -5621 320348 -5615
rect 320108 -5935 320179 -5901
rect 320477 -5935 320547 -5584
rect 320659 -5652 320717 -5646
rect 320659 -5686 320671 -5652
rect 320659 -5692 320717 -5686
rect 320659 -5852 320717 -5846
rect 320659 -5886 320671 -5852
rect 320659 -5892 320717 -5886
rect 320846 -5901 320916 -5514
rect 321198 -5514 321232 -5513
rect 321620 -5513 321655 -5496
rect 321935 -5513 321970 -5496
rect 321620 -5514 321654 -5513
rect 321198 -5550 321268 -5514
rect 321028 -5581 321086 -5575
rect 321028 -5615 321040 -5581
rect 321215 -5584 321286 -5550
rect 321028 -5621 321086 -5615
rect 320846 -5935 320917 -5901
rect 321215 -5935 321285 -5584
rect 321397 -5652 321455 -5646
rect 321397 -5686 321409 -5652
rect 321397 -5692 321455 -5686
rect 321397 -5852 321455 -5846
rect 321397 -5886 321409 -5852
rect 321397 -5892 321455 -5886
rect 321584 -5901 321654 -5514
rect 321936 -5514 321970 -5513
rect 322358 -5514 322393 -5496
rect 321936 -5550 322006 -5514
rect 322322 -5529 322393 -5514
rect 321766 -5581 321824 -5575
rect 321766 -5615 321778 -5581
rect 321953 -5584 322024 -5550
rect 321766 -5621 321824 -5615
rect 321584 -5935 321655 -5901
rect 321953 -5935 322023 -5584
rect 322135 -5652 322193 -5646
rect 322135 -5686 322147 -5652
rect 322135 -5692 322193 -5686
rect 322135 -5852 322193 -5846
rect 322135 -5886 322147 -5852
rect 322135 -5892 322193 -5886
rect 2825 -5971 2882 -5935
rect 2957 -5988 3119 -5954
rect 4012 -5971 4065 -5935
rect 5860 -5971 5913 -5935
rect 7708 -5971 7761 -5935
rect 9556 -5971 9609 -5935
rect 11404 -5971 11457 -5935
rect 13252 -5971 13305 -5935
rect 15100 -5971 15153 -5935
rect 16948 -5971 17001 -5935
rect 18796 -5971 18849 -5935
rect 20644 -5971 20697 -5935
rect 22492 -5971 22545 -5935
rect 24340 -5971 24393 -5935
rect 26188 -5971 26241 -5935
rect 28036 -5971 28089 -5935
rect 29884 -5971 29937 -5935
rect 31732 -5971 31785 -5935
rect 33580 -5971 33633 -5935
rect 35428 -5971 35481 -5935
rect 37276 -5971 37329 -5935
rect 39124 -5971 39177 -5935
rect 40972 -5971 41025 -5935
rect 42820 -5971 42873 -5935
rect 44668 -5971 44721 -5935
rect 46516 -5971 46569 -5935
rect 48364 -5971 48417 -5935
rect 50212 -5971 50265 -5935
rect 52060 -5971 52113 -5935
rect 53908 -5971 53961 -5935
rect 55756 -5971 55809 -5935
rect 57604 -5971 57657 -5935
rect 59452 -5971 59505 -5935
rect 61300 -5971 61353 -5935
rect 63148 -5971 63201 -5935
rect 64996 -5971 65049 -5935
rect 66844 -5971 66897 -5935
rect 68692 -5971 68745 -5935
rect 70540 -5971 70593 -5935
rect 72388 -5971 72441 -5935
rect 74236 -5971 74289 -5935
rect 76084 -5971 76137 -5935
rect 77932 -5971 77985 -5935
rect 79780 -5971 79833 -5935
rect 81628 -5971 81681 -5935
rect 83476 -5971 83529 -5935
rect 85324 -5971 85377 -5935
rect 87172 -5971 87225 -5935
rect 89020 -5971 89073 -5935
rect 90868 -5971 90921 -5935
rect 92716 -5971 92769 -5935
rect 94564 -5971 94617 -5935
rect 96412 -5971 96465 -5935
rect 98260 -5971 98313 -5935
rect 100108 -5971 100161 -5935
rect 101956 -5971 102009 -5935
rect 103804 -5971 103857 -5935
rect 105652 -5971 105705 -5935
rect 107500 -5971 107553 -5935
rect 109348 -5971 109401 -5935
rect 111196 -5971 111249 -5935
rect 113044 -5971 113097 -5935
rect 114892 -5971 114945 -5935
rect 116740 -5971 116793 -5935
rect 118588 -5971 118641 -5935
rect 120436 -5971 120489 -5935
rect 122284 -5971 122337 -5935
rect 124132 -5971 124185 -5935
rect 125980 -5971 126033 -5935
rect 127828 -5971 127881 -5935
rect 129676 -5971 129729 -5935
rect 131524 -5971 131577 -5935
rect 133372 -5971 133425 -5935
rect 135220 -5971 135273 -5935
rect 137068 -5971 137121 -5935
rect 138916 -5971 138969 -5935
rect 140764 -5971 140817 -5935
rect 142612 -5971 142665 -5935
rect 144460 -5971 144513 -5935
rect 146308 -5971 146361 -5935
rect 148156 -5971 148209 -5935
rect 150004 -5971 150057 -5935
rect 151852 -5971 151905 -5935
rect 153700 -5971 153753 -5935
rect 155548 -5971 155601 -5935
rect 157396 -5971 157449 -5935
rect 159244 -5971 159297 -5935
rect 161092 -5971 161145 -5935
rect 162940 -5971 162993 -5935
rect 164788 -5971 164841 -5935
rect 166636 -5971 166689 -5935
rect 168484 -5971 168537 -5935
rect 170332 -5971 170385 -5935
rect 172180 -5971 172233 -5935
rect 174028 -5971 174081 -5935
rect 175876 -5971 175929 -5935
rect 177724 -5971 177777 -5935
rect 179519 -5971 179572 -5935
rect 179888 -5971 179941 -5935
rect 180257 -5971 180310 -5935
rect 180626 -5971 180679 -5935
rect 180995 -5971 181048 -5935
rect 181364 -5971 181417 -5935
rect 181733 -5971 181786 -5935
rect 182102 -5971 182155 -5935
rect 182471 -5971 182524 -5935
rect 182840 -5971 182893 -5935
rect 183209 -5971 183262 -5935
rect 183578 -5971 183631 -5935
rect 183947 -5971 184000 -5935
rect 184316 -5971 184369 -5935
rect 184685 -5971 184738 -5935
rect 185054 -5971 185107 -5935
rect 185423 -5971 185476 -5935
rect 185792 -5971 185845 -5935
rect 186161 -5971 186214 -5935
rect 186530 -5971 186583 -5935
rect 186899 -5971 186952 -5935
rect 187268 -5971 187321 -5935
rect 187637 -5971 187690 -5935
rect 188006 -5971 188059 -5935
rect 188375 -5971 188428 -5935
rect 188744 -5971 188797 -5935
rect 189113 -5971 189166 -5935
rect 189482 -5971 189535 -5935
rect 189851 -5971 189904 -5935
rect 190220 -5971 190273 -5935
rect 190589 -5971 190642 -5935
rect 190958 -5971 191011 -5935
rect 191327 -5971 191380 -5935
rect 191696 -5971 191749 -5935
rect 192065 -5971 192118 -5935
rect 192434 -5971 192487 -5935
rect 192803 -5971 192856 -5935
rect 193172 -5971 193225 -5935
rect 193541 -5971 193594 -5935
rect 193910 -5971 193963 -5935
rect 194279 -5971 194332 -5935
rect 194648 -5971 194701 -5935
rect 195017 -5971 195070 -5935
rect 195386 -5971 195439 -5935
rect 195755 -5971 195808 -5935
rect 196124 -5971 196177 -5935
rect 196493 -5971 196546 -5935
rect 196862 -5971 196915 -5935
rect 197231 -5971 197284 -5935
rect 197600 -5971 197653 -5935
rect 197969 -5971 198022 -5935
rect 198338 -5971 198391 -5935
rect 198707 -5971 198760 -5935
rect 199076 -5971 199129 -5935
rect 199445 -5971 199498 -5935
rect 199814 -5971 199867 -5935
rect 200183 -5971 200236 -5935
rect 200552 -5971 200605 -5935
rect 200921 -5971 200974 -5935
rect 201290 -5971 201343 -5935
rect 201659 -5971 201712 -5935
rect 202028 -5971 202081 -5935
rect 202397 -5971 202450 -5935
rect 202766 -5971 202819 -5935
rect 203135 -5971 203188 -5935
rect 203504 -5971 203557 -5935
rect 203873 -5971 203926 -5935
rect 204242 -5971 204295 -5935
rect 204611 -5971 204664 -5935
rect 204980 -5971 205033 -5935
rect 205349 -5971 205402 -5935
rect 205718 -5971 205771 -5935
rect 206087 -5971 206140 -5935
rect 206456 -5971 206509 -5935
rect 206825 -5971 206878 -5935
rect 207194 -5971 207247 -5935
rect 207563 -5971 207616 -5935
rect 207932 -5971 207985 -5935
rect 208301 -5971 208354 -5935
rect 208670 -5971 208723 -5935
rect 209039 -5971 209092 -5935
rect 209408 -5971 209461 -5935
rect 209777 -5971 209830 -5935
rect 210146 -5971 210199 -5935
rect 210515 -5971 210568 -5935
rect 210884 -5971 210937 -5935
rect 211253 -5971 211306 -5935
rect 211622 -5971 211675 -5935
rect 211991 -5971 212044 -5935
rect 212360 -5971 212413 -5935
rect 212729 -5971 212782 -5935
rect 213098 -5971 213151 -5935
rect 213467 -5971 213520 -5935
rect 213836 -5971 213889 -5935
rect 214205 -5971 214258 -5935
rect 214574 -5971 214627 -5935
rect 214943 -5971 214996 -5935
rect 215312 -5971 215365 -5935
rect 215681 -5971 215734 -5935
rect 216050 -5971 216103 -5935
rect 216419 -5971 216472 -5935
rect 216788 -5971 216841 -5935
rect 217157 -5971 217210 -5935
rect 217526 -5971 217579 -5935
rect 217895 -5971 217948 -5935
rect 218264 -5971 218317 -5935
rect 218633 -5971 218686 -5935
rect 219002 -5971 219055 -5935
rect 219371 -5971 219424 -5935
rect 219740 -5971 219793 -5935
rect 220109 -5971 220162 -5935
rect 220478 -5971 220531 -5935
rect 220847 -5971 220900 -5935
rect 221216 -5971 221269 -5935
rect 221585 -5971 221638 -5935
rect 221954 -5971 222007 -5935
rect 222323 -5971 222376 -5935
rect 222692 -5971 222745 -5935
rect 223061 -5971 223114 -5935
rect 223430 -5971 223483 -5935
rect 223799 -5971 223852 -5935
rect 224168 -5971 224221 -5935
rect 224537 -5971 224590 -5935
rect 224906 -5971 224959 -5935
rect 225275 -5971 225328 -5935
rect 225644 -5971 225697 -5935
rect 226013 -5971 226066 -5935
rect 226382 -5971 226435 -5935
rect 226751 -5971 226804 -5935
rect 227120 -5971 227173 -5935
rect 227489 -5971 227542 -5935
rect 227858 -5971 227911 -5935
rect 228227 -5971 228280 -5935
rect 228596 -5971 228649 -5935
rect 228965 -5971 229018 -5935
rect 229334 -5971 229387 -5935
rect 229703 -5971 229756 -5935
rect 230072 -5971 230125 -5935
rect 230441 -5971 230494 -5935
rect 230810 -5971 230863 -5935
rect 231179 -5971 231232 -5935
rect 231548 -5971 231601 -5935
rect 231917 -5971 231970 -5935
rect 232286 -5971 232339 -5935
rect 232655 -5971 232708 -5935
rect 233024 -5971 233077 -5935
rect 233393 -5971 233446 -5935
rect 233762 -5971 233815 -5935
rect 234131 -5971 234184 -5935
rect 234500 -5971 234553 -5935
rect 234869 -5971 234922 -5935
rect 235238 -5971 235291 -5935
rect 235607 -5971 235660 -5935
rect 235976 -5971 236029 -5935
rect 236345 -5971 236398 -5935
rect 236714 -5971 236767 -5935
rect 237083 -5971 237136 -5935
rect 237452 -5971 237505 -5935
rect 237821 -5971 237874 -5935
rect 238190 -5971 238243 -5935
rect 238559 -5971 238612 -5935
rect 238928 -5971 238981 -5935
rect 239297 -5971 239350 -5935
rect 239666 -5971 239719 -5935
rect 240035 -5971 240088 -5935
rect 240404 -5971 240457 -5935
rect 240773 -5971 240826 -5935
rect 241142 -5971 241195 -5935
rect 241511 -5971 241564 -5935
rect 241880 -5971 241933 -5935
rect 242249 -5971 242302 -5935
rect 242618 -5971 242671 -5935
rect 242987 -5971 243040 -5935
rect 243356 -5971 243409 -5935
rect 243725 -5971 243778 -5935
rect 244094 -5971 244147 -5935
rect 244463 -5971 244516 -5935
rect 244832 -5971 244885 -5935
rect 245201 -5971 245254 -5935
rect 245570 -5971 245623 -5935
rect 245939 -5971 245992 -5935
rect 246308 -5971 246361 -5935
rect 246677 -5971 246730 -5935
rect 247046 -5971 247099 -5935
rect 247415 -5971 247468 -5935
rect 247784 -5971 247837 -5935
rect 248153 -5971 248206 -5935
rect 248522 -5971 248575 -5935
rect 248891 -5971 248944 -5935
rect 249260 -5971 249313 -5935
rect 249629 -5971 249682 -5935
rect 249998 -5971 250051 -5935
rect 250367 -5971 250420 -5935
rect 250736 -5971 250789 -5935
rect 251105 -5971 251158 -5935
rect 251474 -5971 251527 -5935
rect 251843 -5971 251896 -5935
rect 252212 -5971 252265 -5935
rect 252581 -5971 252634 -5935
rect 252950 -5971 253003 -5935
rect 253319 -5971 253372 -5935
rect 253688 -5971 253741 -5935
rect 254057 -5971 254110 -5935
rect 254426 -5971 254479 -5935
rect 254795 -5971 254848 -5935
rect 255164 -5971 255217 -5935
rect 255533 -5971 255586 -5935
rect 255902 -5971 255955 -5935
rect 256271 -5971 256324 -5935
rect 256640 -5971 256693 -5935
rect 257009 -5971 257062 -5935
rect 257378 -5971 257431 -5935
rect 257747 -5971 257800 -5935
rect 258116 -5971 258169 -5935
rect 258485 -5971 258538 -5935
rect 258854 -5971 258907 -5935
rect 259223 -5971 259276 -5935
rect 259592 -5971 259645 -5935
rect 259961 -5971 260014 -5935
rect 260330 -5971 260383 -5935
rect 260699 -5971 260752 -5935
rect 261068 -5971 261121 -5935
rect 261437 -5971 261490 -5935
rect 261806 -5971 261859 -5935
rect 262175 -5971 262228 -5935
rect 262544 -5971 262597 -5935
rect 262913 -5971 262966 -5935
rect 263282 -5971 263335 -5935
rect 263651 -5971 263704 -5935
rect 264020 -5971 264073 -5935
rect 264389 -5971 264442 -5935
rect 264758 -5971 264811 -5935
rect 265127 -5971 265180 -5935
rect 265496 -5971 265549 -5935
rect 265865 -5971 265918 -5935
rect 266234 -5971 266287 -5935
rect 266603 -5971 266656 -5935
rect 266972 -5971 267025 -5935
rect 267341 -5971 267394 -5935
rect 267710 -5971 267763 -5935
rect 268079 -5971 268132 -5935
rect 268448 -5971 268501 -5935
rect 268817 -5971 268870 -5935
rect 269186 -5971 269239 -5935
rect 269555 -5971 269608 -5935
rect 269924 -5971 269977 -5935
rect 270293 -5971 270346 -5935
rect 270662 -5971 270715 -5935
rect 271031 -5971 271084 -5935
rect 271400 -5971 271453 -5935
rect 271769 -5971 271822 -5935
rect 272138 -5971 272191 -5935
rect 272507 -5971 272560 -5935
rect 272876 -5971 272929 -5935
rect 273245 -5971 273298 -5935
rect 273614 -5971 273667 -5935
rect 273983 -5971 274036 -5935
rect 274352 -5971 274405 -5935
rect 274721 -5971 274774 -5935
rect 275090 -5971 275143 -5935
rect 275459 -5971 275512 -5935
rect 275828 -5971 275881 -5935
rect 276197 -5971 276250 -5935
rect 276566 -5971 276619 -5935
rect 276935 -5971 276988 -5935
rect 277304 -5971 277357 -5935
rect 277673 -5971 277726 -5935
rect 278042 -5971 278095 -5935
rect 278411 -5971 278464 -5935
rect 278780 -5971 278833 -5935
rect 279149 -5971 279202 -5935
rect 279518 -5971 279571 -5935
rect 279887 -5971 279940 -5935
rect 280256 -5971 280309 -5935
rect 280625 -5971 280678 -5935
rect 280994 -5971 281047 -5935
rect 281363 -5971 281416 -5935
rect 281732 -5971 281785 -5935
rect 282101 -5971 282154 -5935
rect 282470 -5971 282523 -5935
rect 282839 -5971 282892 -5935
rect 283208 -5971 283261 -5935
rect 283577 -5971 283630 -5935
rect 283946 -5971 283999 -5935
rect 284315 -5971 284368 -5935
rect 284684 -5971 284737 -5935
rect 285053 -5971 285106 -5935
rect 285422 -5971 285475 -5935
rect 285791 -5971 285844 -5935
rect 286160 -5971 286213 -5935
rect 286529 -5971 286582 -5935
rect 286898 -5971 286951 -5935
rect 287267 -5971 287320 -5935
rect 287636 -5971 287689 -5935
rect 288005 -5971 288058 -5935
rect 288374 -5971 288427 -5935
rect 288743 -5971 288796 -5935
rect 289112 -5971 289165 -5935
rect 289481 -5971 289534 -5935
rect 289850 -5971 289903 -5935
rect 290219 -5971 290272 -5935
rect 290588 -5971 290641 -5935
rect 290957 -5971 291010 -5935
rect 291326 -5971 291379 -5935
rect 291695 -5971 291748 -5935
rect 292064 -5971 292117 -5935
rect 292433 -5971 292486 -5935
rect 292802 -5971 292855 -5935
rect 293171 -5971 293224 -5935
rect 293540 -5971 293593 -5935
rect 293909 -5971 293962 -5935
rect 294278 -5971 294331 -5935
rect 294647 -5971 294700 -5935
rect 295016 -5971 295069 -5935
rect 295385 -5971 295438 -5935
rect 295754 -5971 295807 -5935
rect 296123 -5971 296176 -5935
rect 296492 -5971 296545 -5935
rect 296861 -5971 296914 -5935
rect 297230 -5971 297283 -5935
rect 297599 -5971 297652 -5935
rect 297968 -5971 298021 -5935
rect 298337 -5971 298390 -5935
rect 298706 -5971 298759 -5935
rect 299075 -5971 299128 -5935
rect 299444 -5971 299497 -5935
rect 299813 -5971 299866 -5935
rect 300182 -5971 300235 -5935
rect 300551 -5971 300604 -5935
rect 300920 -5971 300973 -5935
rect 301289 -5971 301342 -5935
rect 301658 -5971 301711 -5935
rect 302027 -5971 302080 -5935
rect 302396 -5971 302449 -5935
rect 302765 -5971 302818 -5935
rect 303134 -5971 303187 -5935
rect 303503 -5971 303556 -5935
rect 303872 -5971 303925 -5935
rect 304241 -5971 304294 -5935
rect 304610 -5971 304663 -5935
rect 304979 -5971 305032 -5935
rect 305348 -5971 305401 -5935
rect 305717 -5971 305770 -5935
rect 306086 -5971 306139 -5935
rect 306455 -5971 306508 -5935
rect 306824 -5971 306877 -5935
rect 307193 -5971 307246 -5935
rect 307562 -5971 307615 -5935
rect 307931 -5971 307984 -5935
rect 308300 -5971 308353 -5935
rect 308669 -5971 308722 -5935
rect 309038 -5971 309091 -5935
rect 309407 -5971 309460 -5935
rect 309776 -5971 309829 -5935
rect 310145 -5971 310198 -5935
rect 310514 -5971 310567 -5935
rect 310883 -5971 310936 -5935
rect 311252 -5971 311305 -5935
rect 311621 -5971 311674 -5935
rect 311990 -5971 312043 -5935
rect 312359 -5971 312412 -5935
rect 312728 -5971 312781 -5935
rect 313097 -5971 313150 -5935
rect 313466 -5971 313519 -5935
rect 313835 -5971 313888 -5935
rect 314204 -5971 314257 -5935
rect 314573 -5971 314626 -5935
rect 314942 -5971 314995 -5935
rect 315311 -5971 315364 -5935
rect 315680 -5971 315733 -5935
rect 316049 -5971 316102 -5935
rect 316418 -5971 316471 -5935
rect 316787 -5971 316840 -5935
rect 317156 -5971 317209 -5935
rect 317525 -5971 317578 -5935
rect 317894 -5971 317947 -5935
rect 318263 -5971 318316 -5935
rect 318632 -5971 318685 -5935
rect 319001 -5971 319054 -5935
rect 319370 -5971 319423 -5935
rect 319739 -5971 319792 -5935
rect 320108 -5971 320161 -5935
rect 320477 -5971 320530 -5935
rect 320846 -5971 320899 -5935
rect 321215 -5971 321268 -5935
rect 321584 -5971 321637 -5935
rect 321953 -5971 322006 -5935
rect 322322 -5988 322392 -5529
rect 322504 -5597 322562 -5591
rect 322504 -5631 322516 -5597
rect 322504 -5637 322562 -5631
rect 322674 -5638 322708 -5584
rect 323096 -5635 323131 -5601
rect 322504 -5905 322562 -5899
rect 322504 -5939 322516 -5905
rect 322504 -5945 322562 -5939
rect 322322 -6024 322375 -5988
rect 322693 -6041 322708 -5638
rect 322727 -5672 322762 -5638
rect 322727 -6041 322761 -5672
rect 322873 -5740 322931 -5734
rect 322873 -5774 322885 -5740
rect 322873 -5780 322931 -5774
rect 322873 -5958 322931 -5952
rect 322873 -5992 322885 -5958
rect 322873 -5998 322931 -5992
rect 322727 -6075 322742 -6041
rect 323062 -6094 323077 -5638
rect 323096 -6094 323130 -5635
rect 323242 -5703 323300 -5697
rect 323242 -5737 323254 -5703
rect 323242 -5743 323300 -5737
rect 323412 -5744 323446 -5690
rect 323834 -5741 323869 -5707
rect 323242 -6011 323300 -6005
rect 323242 -6045 323254 -6011
rect 323242 -6051 323300 -6045
rect 323096 -6128 323111 -6094
rect 323431 -6147 323446 -5744
rect 323465 -5778 323500 -5744
rect 323465 -6147 323499 -5778
rect 323611 -5846 323669 -5840
rect 323611 -5880 323623 -5846
rect 323611 -5886 323669 -5880
rect 323611 -6064 323669 -6058
rect 323611 -6098 323623 -6064
rect 323611 -6104 323669 -6098
rect 323465 -6181 323480 -6147
rect 323800 -6200 323815 -5744
rect 323834 -6200 323868 -5741
rect 323980 -5809 324038 -5803
rect 323980 -5843 323992 -5809
rect 323980 -5849 324038 -5843
rect 324150 -5850 324184 -5796
rect 323980 -6117 324038 -6111
rect 323980 -6151 323992 -6117
rect 323980 -6157 324038 -6151
rect 323834 -6234 323849 -6200
rect 324169 -6253 324184 -5850
rect 324203 -5884 324238 -5850
rect 324518 -5884 324553 -5867
rect 324203 -6253 324237 -5884
rect 324519 -5885 324553 -5884
rect 324519 -5921 324589 -5885
rect 324349 -5952 324407 -5946
rect 324349 -5986 324361 -5952
rect 324536 -5955 324607 -5921
rect 324887 -5955 324922 -5921
rect 324349 -5992 324407 -5986
rect 324349 -6170 324407 -6164
rect 324349 -6204 324361 -6170
rect 324349 -6210 324407 -6204
rect 324203 -6287 324218 -6253
rect 324536 -6306 324606 -5955
rect 324888 -5974 324922 -5955
rect 324718 -6023 324776 -6017
rect 324718 -6057 324730 -6023
rect 324718 -6063 324776 -6057
rect 324718 -6223 324776 -6217
rect 324718 -6257 324730 -6223
rect 324718 -6263 324776 -6257
rect 324536 -6342 324589 -6306
rect 324907 -6359 324922 -5974
rect 324941 -6008 324976 -5974
rect 325256 -6008 325291 -5974
rect 324941 -6359 324975 -6008
rect 325257 -6027 325291 -6008
rect 325087 -6076 325145 -6070
rect 325087 -6110 325099 -6076
rect 325087 -6116 325145 -6110
rect 325087 -6276 325145 -6270
rect 325087 -6310 325099 -6276
rect 325087 -6316 325145 -6310
rect 324941 -6393 324956 -6359
rect 325276 -6412 325291 -6027
rect 325310 -6061 325345 -6027
rect 325625 -6061 325660 -6027
rect 325310 -6412 325344 -6061
rect 325626 -6080 325660 -6061
rect 325456 -6129 325514 -6123
rect 325456 -6163 325468 -6129
rect 325456 -6169 325514 -6163
rect 325456 -6329 325514 -6323
rect 325456 -6363 325468 -6329
rect 325456 -6369 325514 -6363
rect 325310 -6446 325325 -6412
rect 325645 -6465 325660 -6080
rect 325679 -6114 325714 -6080
rect 325679 -6465 325713 -6114
rect 325825 -6182 325883 -6176
rect 325825 -6216 325837 -6182
rect 325825 -6222 325883 -6216
rect 325825 -6382 325883 -6376
rect 325825 -6416 325837 -6382
rect 325825 -6422 325883 -6416
rect 325679 -6499 325694 -6465
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use inverter  inverter_0
timestamp 1728247082
transform 1 0 0 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_1
timestamp 1728247082
transform 1 0 1848 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_2
timestamp 1728247082
transform 1 0 3696 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_3
timestamp 1728247082
transform 1 0 5544 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_4
timestamp 1728247082
transform 1 0 7392 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_5
timestamp 1728247082
transform 1 0 9240 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_6
timestamp 1728247082
transform 1 0 11088 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_7
timestamp 1728247082
transform 1 0 12936 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_8
timestamp 1728247082
transform 1 0 14784 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_9
timestamp 1728247082
transform 1 0 16632 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_10
timestamp 1728247082
transform 1 0 18480 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_11
timestamp 1728247082
transform 1 0 20328 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_12
timestamp 1728247082
transform 1 0 22176 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_13
timestamp 1728247082
transform 1 0 24024 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_14
timestamp 1728247082
transform 1 0 25872 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_15
timestamp 1728247082
transform 1 0 27720 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_16
timestamp 1728247082
transform 1 0 29568 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_17
timestamp 1728247082
transform 1 0 31416 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_18
timestamp 1728247082
transform 1 0 33264 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_19
timestamp 1728247082
transform 1 0 35112 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_20
timestamp 1728247082
transform 1 0 36960 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_21
timestamp 1728247082
transform 1 0 38808 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_22
timestamp 1728247082
transform 1 0 40656 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_23
timestamp 1728247082
transform 1 0 42504 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_24
timestamp 1728247082
transform 1 0 44352 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_25
timestamp 1728247082
transform 1 0 46200 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_26
timestamp 1728247082
transform 1 0 48048 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_27
timestamp 1728247082
transform 1 0 49896 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_28
timestamp 1728247082
transform 1 0 51744 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_29
timestamp 1728247082
transform 1 0 53592 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_30
timestamp 1728247082
transform 1 0 55440 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_31
timestamp 1728247082
transform 1 0 57288 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_32
timestamp 1728247082
transform 1 0 59136 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_33
timestamp 1728247082
transform 1 0 60984 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_34
timestamp 1728247082
transform 1 0 62832 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_35
timestamp 1728247082
transform 1 0 64680 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_36
timestamp 1728247082
transform 1 0 66528 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_37
timestamp 1728247082
transform 1 0 68376 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_38
timestamp 1728247082
transform 1 0 70224 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_39
timestamp 1728247082
transform 1 0 72072 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_40
timestamp 1728247082
transform 1 0 73920 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_41
timestamp 1728247082
transform 1 0 75768 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_42
timestamp 1728247082
transform 1 0 77616 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_43
timestamp 1728247082
transform 1 0 79464 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_44
timestamp 1728247082
transform 1 0 81312 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_45
timestamp 1728247082
transform 1 0 83160 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_46
timestamp 1728247082
transform 1 0 85008 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_47
timestamp 1728247082
transform 1 0 86856 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_48
timestamp 1728247082
transform 1 0 88704 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_49
timestamp 1728247082
transform 1 0 90552 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_50
timestamp 1728247082
transform 1 0 92400 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_51
timestamp 1728247082
transform 1 0 94248 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_52
timestamp 1728247082
transform 1 0 96096 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_53
timestamp 1728247082
transform 1 0 97944 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_54
timestamp 1728247082
transform 1 0 99792 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_55
timestamp 1728247082
transform 1 0 101640 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_56
timestamp 1728247082
transform 1 0 103488 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_57
timestamp 1728247082
transform 1 0 105336 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_58
timestamp 1728247082
transform 1 0 107184 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_59
timestamp 1728247082
transform 1 0 109032 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_60
timestamp 1728247082
transform 1 0 110880 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_61
timestamp 1728247082
transform 1 0 112728 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_62
timestamp 1728247082
transform 1 0 114576 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_63
timestamp 1728247082
transform 1 0 116424 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_64
timestamp 1728247082
transform 1 0 118272 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_65
timestamp 1728247082
transform 1 0 120120 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_66
timestamp 1728247082
transform 1 0 121968 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_67
timestamp 1728247082
transform 1 0 123816 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_68
timestamp 1728247082
transform 1 0 125664 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_69
timestamp 1728247082
transform 1 0 127512 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_70
timestamp 1728247082
transform 1 0 129360 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_71
timestamp 1728247082
transform 1 0 131208 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_72
timestamp 1728247082
transform 1 0 133056 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_73
timestamp 1728247082
transform 1 0 134904 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_74
timestamp 1728247082
transform 1 0 136752 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_75
timestamp 1728247082
transform 1 0 138600 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_76
timestamp 1728247082
transform 1 0 140448 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_77
timestamp 1728247082
transform 1 0 142296 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_78
timestamp 1728247082
transform 1 0 144144 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_79
timestamp 1728247082
transform 1 0 145992 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_80
timestamp 1728247082
transform 1 0 147840 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_81
timestamp 1728247082
transform 1 0 149688 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_82
timestamp 1728247082
transform 1 0 151536 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_83
timestamp 1728247082
transform 1 0 153384 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_84
timestamp 1728247082
transform 1 0 155232 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_85
timestamp 1728247082
transform 1 0 157080 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_86
timestamp 1728247082
transform 1 0 158928 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_87
timestamp 1728247082
transform 1 0 160776 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_88
timestamp 1728247082
transform 1 0 162624 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_89
timestamp 1728247082
transform 1 0 164472 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_90
timestamp 1728247082
transform 1 0 166320 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_91
timestamp 1728247082
transform 1 0 168168 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_92
timestamp 1728247082
transform 1 0 170016 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_93
timestamp 1728247082
transform 1 0 171864 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_94
timestamp 1728247082
transform 1 0 173712 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_95
timestamp 1728247082
transform 1 0 175560 0 1 -4718
box -53 -1306 1795 200
use inverter  inverter_96
timestamp 1728247082
transform 1 0 177408 0 1 -4718
box -53 -1306 1795 200
use passGate_hvt  passGate_hvt_0
timestamp 1728244868
transform 1 0 179203 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_1
timestamp 1728244868
transform 1 0 179941 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_2
timestamp 1728244868
transform 1 0 180679 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_3
timestamp 1728244868
transform 1 0 181417 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_4
timestamp 1728244868
transform 1 0 182155 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_5
timestamp 1728244868
transform 1 0 182893 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_6
timestamp 1728244868
transform 1 0 183631 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_7
timestamp 1728244868
transform 1 0 184369 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_8
timestamp 1728244868
transform 1 0 185107 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_9
timestamp 1728244868
transform 1 0 185845 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_10
timestamp 1728244868
transform 1 0 186583 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_11
timestamp 1728244868
transform 1 0 187321 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_12
timestamp 1728244868
transform 1 0 188059 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_13
timestamp 1728244868
transform 1 0 188797 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_14
timestamp 1728244868
transform 1 0 189535 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_15
timestamp 1728244868
transform 1 0 190273 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_16
timestamp 1728244868
transform 1 0 191011 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_17
timestamp 1728244868
transform 1 0 191749 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_18
timestamp 1728244868
transform 1 0 192487 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_19
timestamp 1728244868
transform 1 0 193225 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_20
timestamp 1728244868
transform 1 0 193963 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_21
timestamp 1728244868
transform 1 0 194701 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_22
timestamp 1728244868
transform 1 0 195439 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_23
timestamp 1728244868
transform 1 0 196177 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_24
timestamp 1728244868
transform 1 0 196915 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_25
timestamp 1728244868
transform 1 0 197653 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_26
timestamp 1728244868
transform 1 0 198391 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_27
timestamp 1728244868
transform 1 0 199129 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_28
timestamp 1728244868
transform 1 0 199867 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_29
timestamp 1728244868
transform 1 0 200605 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_30
timestamp 1728244868
transform 1 0 201343 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_31
timestamp 1728244868
transform 1 0 202081 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_32
timestamp 1728244868
transform 1 0 202819 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_33
timestamp 1728244868
transform 1 0 203557 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_34
timestamp 1728244868
transform 1 0 204295 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_35
timestamp 1728244868
transform 1 0 205033 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_36
timestamp 1728244868
transform 1 0 205771 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_37
timestamp 1728244868
transform 1 0 206509 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_38
timestamp 1728244868
transform 1 0 207247 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_39
timestamp 1728244868
transform 1 0 207985 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_40
timestamp 1728244868
transform 1 0 208723 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_41
timestamp 1728244868
transform 1 0 209461 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_42
timestamp 1728244868
transform 1 0 210199 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_43
timestamp 1728244868
transform 1 0 210937 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_44
timestamp 1728244868
transform 1 0 211675 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_45
timestamp 1728244868
transform 1 0 212413 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_46
timestamp 1728244868
transform 1 0 213151 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_47
timestamp 1728244868
transform 1 0 213889 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_48
timestamp 1728244868
transform 1 0 214627 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_49
timestamp 1728244868
transform 1 0 215365 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_50
timestamp 1728244868
transform 1 0 216103 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_51
timestamp 1728244868
transform 1 0 216841 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_52
timestamp 1728244868
transform 1 0 217579 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_53
timestamp 1728244868
transform 1 0 218317 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_54
timestamp 1728244868
transform 1 0 219055 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_55
timestamp 1728244868
transform 1 0 219793 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_56
timestamp 1728244868
transform 1 0 220531 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_57
timestamp 1728244868
transform 1 0 221269 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_58
timestamp 1728244868
transform 1 0 222007 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_59
timestamp 1728244868
transform 1 0 222745 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_60
timestamp 1728244868
transform 1 0 223483 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_61
timestamp 1728244868
transform 1 0 224221 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_62
timestamp 1728244868
transform 1 0 224959 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_63
timestamp 1728244868
transform 1 0 225697 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_64
timestamp 1728244868
transform 1 0 226435 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_65
timestamp 1728244868
transform 1 0 227173 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_66
timestamp 1728244868
transform 1 0 227911 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_67
timestamp 1728244868
transform 1 0 228649 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_68
timestamp 1728244868
transform 1 0 229387 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_69
timestamp 1728244868
transform 1 0 230125 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_70
timestamp 1728244868
transform 1 0 230863 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_71
timestamp 1728244868
transform 1 0 231601 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_72
timestamp 1728244868
transform 1 0 232339 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_73
timestamp 1728244868
transform 1 0 233077 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_74
timestamp 1728244868
transform 1 0 233815 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_75
timestamp 1728244868
transform 1 0 234553 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_76
timestamp 1728244868
transform 1 0 235291 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_77
timestamp 1728244868
transform 1 0 236029 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_78
timestamp 1728244868
transform 1 0 236767 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_79
timestamp 1728244868
transform 1 0 237505 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_80
timestamp 1728244868
transform 1 0 238243 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_81
timestamp 1728244868
transform 1 0 238981 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_82
timestamp 1728244868
transform 1 0 239719 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_83
timestamp 1728244868
transform 1 0 240457 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_84
timestamp 1728244868
transform 1 0 241195 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_85
timestamp 1728244868
transform 1 0 241933 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_86
timestamp 1728244868
transform 1 0 242671 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_87
timestamp 1728244868
transform 1 0 243409 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_88
timestamp 1728244868
transform 1 0 244147 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_89
timestamp 1728244868
transform 1 0 244885 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_90
timestamp 1728244868
transform 1 0 245623 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_91
timestamp 1728244868
transform 1 0 246361 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_92
timestamp 1728244868
transform 1 0 247099 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_93
timestamp 1728244868
transform 1 0 247837 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_94
timestamp 1728244868
transform 1 0 248575 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_95
timestamp 1728244868
transform 1 0 249313 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_96
timestamp 1728244868
transform 1 0 250051 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_97
timestamp 1728244868
transform 1 0 250789 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_98
timestamp 1728244868
transform 1 0 251527 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_99
timestamp 1728244868
transform 1 0 252265 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_100
timestamp 1728244868
transform 1 0 253003 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_101
timestamp 1728244868
transform 1 0 253741 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_102
timestamp 1728244868
transform 1 0 254479 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_103
timestamp 1728244868
transform 1 0 255217 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_104
timestamp 1728244868
transform 1 0 255955 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_105
timestamp 1728244868
transform 1 0 256693 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_106
timestamp 1728244868
transform 1 0 257431 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_107
timestamp 1728244868
transform 1 0 258169 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_108
timestamp 1728244868
transform 1 0 258907 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_109
timestamp 1728244868
transform 1 0 259645 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_110
timestamp 1728244868
transform 1 0 260383 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_111
timestamp 1728244868
transform 1 0 261121 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_112
timestamp 1728244868
transform 1 0 261859 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_113
timestamp 1728244868
transform 1 0 262597 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_114
timestamp 1728244868
transform 1 0 263335 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_115
timestamp 1728244868
transform 1 0 264073 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_116
timestamp 1728244868
transform 1 0 264811 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_117
timestamp 1728244868
transform 1 0 265549 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_118
timestamp 1728244868
transform 1 0 266287 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_119
timestamp 1728244868
transform 1 0 267025 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_120
timestamp 1728244868
transform 1 0 267763 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_121
timestamp 1728244868
transform 1 0 268501 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_122
timestamp 1728244868
transform 1 0 269239 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_123
timestamp 1728244868
transform 1 0 269977 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_124
timestamp 1728244868
transform 1 0 270715 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_125
timestamp 1728244868
transform 1 0 271453 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_126
timestamp 1728244868
transform 1 0 272191 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_127
timestamp 1728244868
transform 1 0 272929 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_128
timestamp 1728244868
transform 1 0 273667 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_129
timestamp 1728244868
transform 1 0 274405 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_130
timestamp 1728244868
transform 1 0 275143 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_131
timestamp 1728244868
transform 1 0 275881 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_132
timestamp 1728244868
transform 1 0 276619 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_133
timestamp 1728244868
transform 1 0 277357 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_134
timestamp 1728244868
transform 1 0 278095 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_135
timestamp 1728244868
transform 1 0 278833 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_136
timestamp 1728244868
transform 1 0 279571 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_137
timestamp 1728244868
transform 1 0 280309 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_138
timestamp 1728244868
transform 1 0 281047 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_139
timestamp 1728244868
transform 1 0 281785 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_140
timestamp 1728244868
transform 1 0 282523 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_141
timestamp 1728244868
transform 1 0 283261 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_142
timestamp 1728244868
transform 1 0 283999 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_143
timestamp 1728244868
transform 1 0 284737 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_144
timestamp 1728244868
transform 1 0 285475 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_145
timestamp 1728244868
transform 1 0 286213 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_146
timestamp 1728244868
transform 1 0 286951 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_147
timestamp 1728244868
transform 1 0 287689 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_148
timestamp 1728244868
transform 1 0 288427 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_149
timestamp 1728244868
transform 1 0 289165 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_150
timestamp 1728244868
transform 1 0 289903 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_151
timestamp 1728244868
transform 1 0 290641 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_152
timestamp 1728244868
transform 1 0 291379 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_153
timestamp 1728244868
transform 1 0 292117 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_154
timestamp 1728244868
transform 1 0 292855 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_155
timestamp 1728244868
transform 1 0 293593 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_156
timestamp 1728244868
transform 1 0 294331 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_157
timestamp 1728244868
transform 1 0 295069 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_158
timestamp 1728244868
transform 1 0 295807 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_159
timestamp 1728244868
transform 1 0 296545 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_160
timestamp 1728244868
transform 1 0 297283 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_161
timestamp 1728244868
transform 1 0 298021 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_162
timestamp 1728244868
transform 1 0 298759 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_163
timestamp 1728244868
transform 1 0 299497 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_164
timestamp 1728244868
transform 1 0 300235 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_165
timestamp 1728244868
transform 1 0 300973 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_166
timestamp 1728244868
transform 1 0 301711 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_167
timestamp 1728244868
transform 1 0 302449 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_168
timestamp 1728244868
transform 1 0 303187 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_169
timestamp 1728244868
transform 1 0 303925 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_170
timestamp 1728244868
transform 1 0 304663 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_171
timestamp 1728244868
transform 1 0 305401 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_172
timestamp 1728244868
transform 1 0 306139 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_173
timestamp 1728244868
transform 1 0 306877 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_174
timestamp 1728244868
transform 1 0 307615 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_175
timestamp 1728244868
transform 1 0 308353 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_176
timestamp 1728244868
transform 1 0 309091 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_177
timestamp 1728244868
transform 1 0 309829 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_178
timestamp 1728244868
transform 1 0 310567 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_179
timestamp 1728244868
transform 1 0 311305 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_180
timestamp 1728244868
transform 1 0 312043 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_181
timestamp 1728244868
transform 1 0 312781 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_182
timestamp 1728244868
transform 1 0 313519 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_183
timestamp 1728244868
transform 1 0 314257 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_184
timestamp 1728244868
transform 1 0 314995 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_185
timestamp 1728244868
transform 1 0 315733 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_186
timestamp 1728244868
transform 1 0 316471 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_187
timestamp 1728244868
transform 1 0 317209 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_188
timestamp 1728244868
transform 1 0 317947 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_189
timestamp 1728244868
transform 1 0 318685 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_190
timestamp 1728244868
transform 1 0 319423 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_191
timestamp 1728244868
transform 1 0 320161 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_192
timestamp 1728244868
transform 1 0 320899 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  passGate_hvt_193
timestamp 1728244868
transform 1 0 321637 0 1 -3918
box -53 -2106 738 200
use inverter  x1[1]
timestamp 1728247082
transform 1 0 0 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[2]
timestamp 1728247082
transform 1 0 1 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[3]
timestamp 1728247082
transform 1 0 2 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[4]
timestamp 1728247082
transform 1 0 3 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[5]
timestamp 1728247082
transform 1 0 4 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[6]
timestamp 1728247082
transform 1 0 5 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[7]
timestamp 1728247082
transform 1 0 6 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[8]
timestamp 1728247082
transform 1 0 7 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[9]
timestamp 1728247082
transform 1 0 8 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[10]
timestamp 1728247082
transform 1 0 9 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[11]
timestamp 1728247082
transform 1 0 10 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[12]
timestamp 1728247082
transform 1 0 11 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[13]
timestamp 1728247082
transform 1 0 12 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[14]
timestamp 1728247082
transform 1 0 13 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[15]
timestamp 1728247082
transform 1 0 14 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[16]
timestamp 1728247082
transform 1 0 15 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[17]
timestamp 1728247082
transform 1 0 16 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[18]
timestamp 1728247082
transform 1 0 17 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[19]
timestamp 1728247082
transform 1 0 18 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[20]
timestamp 1728247082
transform 1 0 19 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[21]
timestamp 1728247082
transform 1 0 20 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[22]
timestamp 1728247082
transform 1 0 21 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[23]
timestamp 1728247082
transform 1 0 22 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[24]
timestamp 1728247082
transform 1 0 23 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[25]
timestamp 1728247082
transform 1 0 24 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[26]
timestamp 1728247082
transform 1 0 25 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[27]
timestamp 1728247082
transform 1 0 26 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[28]
timestamp 1728247082
transform 1 0 27 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[29]
timestamp 1728247082
transform 1 0 28 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[30]
timestamp 1728247082
transform 1 0 29 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[31]
timestamp 1728247082
transform 1 0 30 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[32]
timestamp 1728247082
transform 1 0 31 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[33]
timestamp 1728247082
transform 1 0 32 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[34]
timestamp 1728247082
transform 1 0 33 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[35]
timestamp 1728247082
transform 1 0 34 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[36]
timestamp 1728247082
transform 1 0 35 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[37]
timestamp 1728247082
transform 1 0 36 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[38]
timestamp 1728247082
transform 1 0 37 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[39]
timestamp 1728247082
transform 1 0 38 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[40]
timestamp 1728247082
transform 1 0 39 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[41]
timestamp 1728247082
transform 1 0 40 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[42]
timestamp 1728247082
transform 1 0 41 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[43]
timestamp 1728247082
transform 1 0 42 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[44]
timestamp 1728247082
transform 1 0 43 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[45]
timestamp 1728247082
transform 1 0 44 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[46]
timestamp 1728247082
transform 1 0 45 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[47]
timestamp 1728247082
transform 1 0 46 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[48]
timestamp 1728247082
transform 1 0 47 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[49]
timestamp 1728247082
transform 1 0 48 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[50]
timestamp 1728247082
transform 1 0 49 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[51]
timestamp 1728247082
transform 1 0 50 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[52]
timestamp 1728247082
transform 1 0 51 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[53]
timestamp 1728247082
transform 1 0 52 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[54]
timestamp 1728247082
transform 1 0 53 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[55]
timestamp 1728247082
transform 1 0 54 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[56]
timestamp 1728247082
transform 1 0 55 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[57]
timestamp 1728247082
transform 1 0 56 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[58]
timestamp 1728247082
transform 1 0 57 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[59]
timestamp 1728247082
transform 1 0 58 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[60]
timestamp 1728247082
transform 1 0 59 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[61]
timestamp 1728247082
transform 1 0 60 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[62]
timestamp 1728247082
transform 1 0 61 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[63]
timestamp 1728247082
transform 1 0 62 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[64]
timestamp 1728247082
transform 1 0 63 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[65]
timestamp 1728247082
transform 1 0 64 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[66]
timestamp 1728247082
transform 1 0 65 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[67]
timestamp 1728247082
transform 1 0 66 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[68]
timestamp 1728247082
transform 1 0 67 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[69]
timestamp 1728247082
transform 1 0 68 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[70]
timestamp 1728247082
transform 1 0 69 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[71]
timestamp 1728247082
transform 1 0 70 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[72]
timestamp 1728247082
transform 1 0 71 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[73]
timestamp 1728247082
transform 1 0 72 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[74]
timestamp 1728247082
transform 1 0 73 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[75]
timestamp 1728247082
transform 1 0 74 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[76]
timestamp 1728247082
transform 1 0 75 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[77]
timestamp 1728247082
transform 1 0 76 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[78]
timestamp 1728247082
transform 1 0 77 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[79]
timestamp 1728247082
transform 1 0 78 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[80]
timestamp 1728247082
transform 1 0 79 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[81]
timestamp 1728247082
transform 1 0 80 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[82]
timestamp 1728247082
transform 1 0 81 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[83]
timestamp 1728247082
transform 1 0 82 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[84]
timestamp 1728247082
transform 1 0 83 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[85]
timestamp 1728247082
transform 1 0 84 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[86]
timestamp 1728247082
transform 1 0 85 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[87]
timestamp 1728247082
transform 1 0 86 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[88]
timestamp 1728247082
transform 1 0 87 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[89]
timestamp 1728247082
transform 1 0 88 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[90]
timestamp 1728247082
transform 1 0 89 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[91]
timestamp 1728247082
transform 1 0 90 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[92]
timestamp 1728247082
transform 1 0 91 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[93]
timestamp 1728247082
transform 1 0 92 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[94]
timestamp 1728247082
transform 1 0 93 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[95]
timestamp 1728247082
transform 1 0 94 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[96]
timestamp 1728247082
transform 1 0 95 0 1 -3600
box -53 -1306 1795 200
use inverter  x1[97]
timestamp 1728247082
transform 1 0 96 0 1 -3600
box -53 -1306 1795 200
use passGate_hvt  x1
timestamp 1728244868
transform 1 0 1769 0 1 -3812
box -53 -2106 738 200
use passGate_hvt  x2
timestamp 1728244868
transform 1 0 1770 0 1 -3812
box -53 -2106 738 200
use passGate_hvt  x2[1]
timestamp 1728244868
transform 1 0 97 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[2]
timestamp 1728244868
transform 1 0 98 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[3]
timestamp 1728244868
transform 1 0 99 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[4]
timestamp 1728244868
transform 1 0 100 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[5]
timestamp 1728244868
transform 1 0 101 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[6]
timestamp 1728244868
transform 1 0 102 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[7]
timestamp 1728244868
transform 1 0 103 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[8]
timestamp 1728244868
transform 1 0 104 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[9]
timestamp 1728244868
transform 1 0 105 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[10]
timestamp 1728244868
transform 1 0 106 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[11]
timestamp 1728244868
transform 1 0 107 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[12]
timestamp 1728244868
transform 1 0 108 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[13]
timestamp 1728244868
transform 1 0 109 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[14]
timestamp 1728244868
transform 1 0 110 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[15]
timestamp 1728244868
transform 1 0 111 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[16]
timestamp 1728244868
transform 1 0 112 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[17]
timestamp 1728244868
transform 1 0 113 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[18]
timestamp 1728244868
transform 1 0 114 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[19]
timestamp 1728244868
transform 1 0 115 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[20]
timestamp 1728244868
transform 1 0 116 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[21]
timestamp 1728244868
transform 1 0 117 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[22]
timestamp 1728244868
transform 1 0 118 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[23]
timestamp 1728244868
transform 1 0 119 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[24]
timestamp 1728244868
transform 1 0 120 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[25]
timestamp 1728244868
transform 1 0 121 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[26]
timestamp 1728244868
transform 1 0 122 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[27]
timestamp 1728244868
transform 1 0 123 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[28]
timestamp 1728244868
transform 1 0 124 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[29]
timestamp 1728244868
transform 1 0 125 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[30]
timestamp 1728244868
transform 1 0 126 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[31]
timestamp 1728244868
transform 1 0 127 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[32]
timestamp 1728244868
transform 1 0 128 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[33]
timestamp 1728244868
transform 1 0 129 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[34]
timestamp 1728244868
transform 1 0 130 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[35]
timestamp 1728244868
transform 1 0 131 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[36]
timestamp 1728244868
transform 1 0 132 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[37]
timestamp 1728244868
transform 1 0 133 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[38]
timestamp 1728244868
transform 1 0 134 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[39]
timestamp 1728244868
transform 1 0 135 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[40]
timestamp 1728244868
transform 1 0 136 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[41]
timestamp 1728244868
transform 1 0 137 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[42]
timestamp 1728244868
transform 1 0 138 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[43]
timestamp 1728244868
transform 1 0 139 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[44]
timestamp 1728244868
transform 1 0 140 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[45]
timestamp 1728244868
transform 1 0 141 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[46]
timestamp 1728244868
transform 1 0 142 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[47]
timestamp 1728244868
transform 1 0 143 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[48]
timestamp 1728244868
transform 1 0 144 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[49]
timestamp 1728244868
transform 1 0 145 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[50]
timestamp 1728244868
transform 1 0 146 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[51]
timestamp 1728244868
transform 1 0 147 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[52]
timestamp 1728244868
transform 1 0 148 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[53]
timestamp 1728244868
transform 1 0 149 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[54]
timestamp 1728244868
transform 1 0 150 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[55]
timestamp 1728244868
transform 1 0 151 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[56]
timestamp 1728244868
transform 1 0 152 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[57]
timestamp 1728244868
transform 1 0 153 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[58]
timestamp 1728244868
transform 1 0 154 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[59]
timestamp 1728244868
transform 1 0 155 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[60]
timestamp 1728244868
transform 1 0 156 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[61]
timestamp 1728244868
transform 1 0 157 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[62]
timestamp 1728244868
transform 1 0 158 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[63]
timestamp 1728244868
transform 1 0 159 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[64]
timestamp 1728244868
transform 1 0 160 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[65]
timestamp 1728244868
transform 1 0 161 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[66]
timestamp 1728244868
transform 1 0 162 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[67]
timestamp 1728244868
transform 1 0 163 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[68]
timestamp 1728244868
transform 1 0 164 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[69]
timestamp 1728244868
transform 1 0 165 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[70]
timestamp 1728244868
transform 1 0 166 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[71]
timestamp 1728244868
transform 1 0 167 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[72]
timestamp 1728244868
transform 1 0 168 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[73]
timestamp 1728244868
transform 1 0 169 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[74]
timestamp 1728244868
transform 1 0 170 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[75]
timestamp 1728244868
transform 1 0 171 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[76]
timestamp 1728244868
transform 1 0 172 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[77]
timestamp 1728244868
transform 1 0 173 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[78]
timestamp 1728244868
transform 1 0 174 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[79]
timestamp 1728244868
transform 1 0 175 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[80]
timestamp 1728244868
transform 1 0 176 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[81]
timestamp 1728244868
transform 1 0 177 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[82]
timestamp 1728244868
transform 1 0 178 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[83]
timestamp 1728244868
transform 1 0 179 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[84]
timestamp 1728244868
transform 1 0 180 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[85]
timestamp 1728244868
transform 1 0 181 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[86]
timestamp 1728244868
transform 1 0 182 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[87]
timestamp 1728244868
transform 1 0 183 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[88]
timestamp 1728244868
transform 1 0 184 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[89]
timestamp 1728244868
transform 1 0 185 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[90]
timestamp 1728244868
transform 1 0 186 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[91]
timestamp 1728244868
transform 1 0 187 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[92]
timestamp 1728244868
transform 1 0 188 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[93]
timestamp 1728244868
transform 1 0 189 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[94]
timestamp 1728244868
transform 1 0 190 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[95]
timestamp 1728244868
transform 1 0 191 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[96]
timestamp 1728244868
transform 1 0 192 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x2[97]
timestamp 1728244868
transform 1 0 193 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3
timestamp 1728244868
transform 1 0 2509 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  x3[1]
timestamp 1728244868
transform 1 0 194 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[2]
timestamp 1728244868
transform 1 0 195 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[3]
timestamp 1728244868
transform 1 0 196 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[4]
timestamp 1728244868
transform 1 0 197 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[5]
timestamp 1728244868
transform 1 0 198 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[6]
timestamp 1728244868
transform 1 0 199 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[7]
timestamp 1728244868
transform 1 0 200 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[8]
timestamp 1728244868
transform 1 0 201 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[9]
timestamp 1728244868
transform 1 0 202 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[10]
timestamp 1728244868
transform 1 0 203 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[11]
timestamp 1728244868
transform 1 0 204 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[12]
timestamp 1728244868
transform 1 0 205 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[13]
timestamp 1728244868
transform 1 0 206 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[14]
timestamp 1728244868
transform 1 0 207 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[15]
timestamp 1728244868
transform 1 0 208 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[16]
timestamp 1728244868
transform 1 0 209 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[17]
timestamp 1728244868
transform 1 0 210 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[18]
timestamp 1728244868
transform 1 0 211 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[19]
timestamp 1728244868
transform 1 0 212 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[20]
timestamp 1728244868
transform 1 0 213 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[21]
timestamp 1728244868
transform 1 0 214 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[22]
timestamp 1728244868
transform 1 0 215 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[23]
timestamp 1728244868
transform 1 0 216 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[24]
timestamp 1728244868
transform 1 0 217 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[25]
timestamp 1728244868
transform 1 0 218 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[26]
timestamp 1728244868
transform 1 0 219 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[27]
timestamp 1728244868
transform 1 0 220 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[28]
timestamp 1728244868
transform 1 0 221 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[29]
timestamp 1728244868
transform 1 0 222 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[30]
timestamp 1728244868
transform 1 0 223 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[31]
timestamp 1728244868
transform 1 0 224 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[32]
timestamp 1728244868
transform 1 0 225 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[33]
timestamp 1728244868
transform 1 0 226 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[34]
timestamp 1728244868
transform 1 0 227 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[35]
timestamp 1728244868
transform 1 0 228 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[36]
timestamp 1728244868
transform 1 0 229 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[37]
timestamp 1728244868
transform 1 0 230 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[38]
timestamp 1728244868
transform 1 0 231 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[39]
timestamp 1728244868
transform 1 0 232 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[40]
timestamp 1728244868
transform 1 0 233 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[41]
timestamp 1728244868
transform 1 0 234 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[42]
timestamp 1728244868
transform 1 0 235 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[43]
timestamp 1728244868
transform 1 0 236 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[44]
timestamp 1728244868
transform 1 0 237 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[45]
timestamp 1728244868
transform 1 0 238 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[46]
timestamp 1728244868
transform 1 0 239 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[47]
timestamp 1728244868
transform 1 0 240 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[48]
timestamp 1728244868
transform 1 0 241 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[49]
timestamp 1728244868
transform 1 0 242 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[50]
timestamp 1728244868
transform 1 0 243 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[51]
timestamp 1728244868
transform 1 0 244 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[52]
timestamp 1728244868
transform 1 0 245 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[53]
timestamp 1728244868
transform 1 0 246 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[54]
timestamp 1728244868
transform 1 0 247 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[55]
timestamp 1728244868
transform 1 0 248 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[56]
timestamp 1728244868
transform 1 0 249 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[57]
timestamp 1728244868
transform 1 0 250 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[58]
timestamp 1728244868
transform 1 0 251 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[59]
timestamp 1728244868
transform 1 0 252 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[60]
timestamp 1728244868
transform 1 0 253 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[61]
timestamp 1728244868
transform 1 0 254 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[62]
timestamp 1728244868
transform 1 0 255 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[63]
timestamp 1728244868
transform 1 0 256 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[64]
timestamp 1728244868
transform 1 0 257 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[65]
timestamp 1728244868
transform 1 0 258 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[66]
timestamp 1728244868
transform 1 0 259 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[67]
timestamp 1728244868
transform 1 0 260 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[68]
timestamp 1728244868
transform 1 0 261 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[69]
timestamp 1728244868
transform 1 0 262 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[70]
timestamp 1728244868
transform 1 0 263 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[71]
timestamp 1728244868
transform 1 0 264 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[72]
timestamp 1728244868
transform 1 0 265 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[73]
timestamp 1728244868
transform 1 0 266 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[74]
timestamp 1728244868
transform 1 0 267 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[75]
timestamp 1728244868
transform 1 0 268 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[76]
timestamp 1728244868
transform 1 0 269 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[77]
timestamp 1728244868
transform 1 0 270 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[78]
timestamp 1728244868
transform 1 0 271 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[79]
timestamp 1728244868
transform 1 0 272 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[80]
timestamp 1728244868
transform 1 0 273 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[81]
timestamp 1728244868
transform 1 0 274 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[82]
timestamp 1728244868
transform 1 0 275 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[83]
timestamp 1728244868
transform 1 0 276 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[84]
timestamp 1728244868
transform 1 0 277 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[85]
timestamp 1728244868
transform 1 0 278 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[86]
timestamp 1728244868
transform 1 0 279 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[87]
timestamp 1728244868
transform 1 0 280 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[88]
timestamp 1728244868
transform 1 0 281 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[89]
timestamp 1728244868
transform 1 0 282 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[90]
timestamp 1728244868
transform 1 0 283 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[91]
timestamp 1728244868
transform 1 0 284 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[92]
timestamp 1728244868
transform 1 0 285 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[93]
timestamp 1728244868
transform 1 0 286 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[94]
timestamp 1728244868
transform 1 0 287 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[95]
timestamp 1728244868
transform 1 0 288 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[96]
timestamp 1728244868
transform 1 0 289 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x3[97]
timestamp 1728244868
transform 1 0 290 0 1 -3600
box -53 -2106 738 200
use passGate_hvt  x4
timestamp 1728244868
transform 1 0 1029 0 1 -3706
box -53 -2106 738 200
use passGate_hvt  x5
timestamp 1728244868
transform 1 0 1030 0 1 -3706
box -53 -2106 738 200
use passGate_hvt  x6
timestamp 1728244868
transform 1 0 2510 0 1 -3918
box -53 -2106 738 200
use inverter  x7
timestamp 1728247082
transform 1 0 2511 0 1 -3918
box -53 -1306 1795 200
use passGate_hvt  x8
timestamp 1728244868
transform 1 0 2512 0 1 -3918
box -53 -2106 738 200
use passGate_hvt  x9
timestamp 1728244868
transform 1 0 2513 0 1 -3918
box -53 -2106 738 200
use sky130_fd_pr__nfet_01v8_4A3DHF  XM1
timestamp 0
transform 1 0 324747 0 1 -6140
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_4A3DHF  XM2
timestamp 0
transform 1 0 325116 0 1 -6193
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_hvt_HVTLRR  XM3
timestamp 0
transform 1 0 322533 0 1 -5768
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_hvt_SNMNDE  XM4
timestamp 0
transform 1 0 322902 0 1 -5866
box -211 -264 211 264
use sky130_fd_pr__nfet_01v8_4A3DHF  XM5
timestamp 0
transform 1 0 325485 0 1 -6246
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_4A3DHF  XM6
timestamp 0
transform 1 0 325854 0 1 -6299
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_hvt_HVTLRR  XM7
timestamp 0
transform 1 0 323271 0 1 -5874
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_hvt_SNMNDE  XM8
timestamp 0
transform 1 0 323640 0 1 -5972
box -211 -264 211 264
use sky130_fd_pr__nfet_01v8_4A3DHF  XM9
timestamp 0
transform 1 0 326223 0 1 -6352
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_hvt_HVTLRR  XM10
timestamp 0
transform 1 0 324009 0 1 -5980
box -211 -309 211 309
use sky130_fd_pr__pfet_01v8_hvt_SNMNDE  XM11
timestamp 0
transform 1 0 324378 0 1 -6078
box -211 -264 211 264
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 DUT_FOOTER
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 DUT_HEADER
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 DUT_GATE
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 NOT_RO_CON
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 RO_CON
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 DRAIN_SENSE
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 {A\[1\]}
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 DRAIN_FORCE
port 9 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 {A\[1\]}
<< end >>
