magic
tech sky130
timestamp 1729529908
<< checkpaint >>
<< l68d20 >>
<< l69d20 >>
<< l68d44 >>
<< end >>
