* Extracted by KLayout with SKY130 LVS runset on : 10/11/2024 16:01

.SUBCKT RO_LVT_13St_x10 RON GND DUT_Gate RO DUT_Header DUT_Footer Drain_Force
+ VDD Drain_Sense OUT
M$1 \$29 \$23 \$16 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$5 VDD RON \$29 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$45 \$30 \$16 \$18 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$49 VDD DUT_Footer \$30 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$89 \$18 RO Drain_Sense VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$93 \$18 RO Drain_Force VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$97 \$32 \$18 \$19 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$101 VDD RON \$32 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$141 \$78 VDD \$23 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$142 \$79 VDD \$23 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$143 VDD \$69 \$23 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$147 \$80 VDD \$69 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$148 \$81 VDD \$69 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$149 VDD \$70 \$69 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$153 \$82 VDD \$70 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$154 \$83 VDD \$70 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$155 VDD \$71 \$70 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$159 \$16 RO DUT_Gate VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$160 \$84 VDD \$71 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$161 \$16 RO \$17 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$162 \$85 VDD \$71 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$163 VDD \$72 \$71 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$167 \$86 VDD \$72 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$168 \$87 VDD \$72 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$169 VDD \$73 \$72 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$173 \$88 VDD \$73 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$174 \$89 VDD \$73 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$175 VDD \$74 \$73 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$179 \$90 VDD \$74 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$180 \$91 VDD \$74 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$181 VDD \$75 \$74 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$185 \$92 VDD \$75 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$186 \$93 VDD \$75 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$187 VDD \$76 \$75 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$191 \$94 VDD \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$192 \$95 VDD \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$193 VDD OUT \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$197 \$96 VDD OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$198 \$97 VDD OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$199 VDD \$19 OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$203 \$19 VDD GND VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$204 \$19 VDD \$20 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$205 \$16 \$23 \$4 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.533e+12 AD=1.533e+12 PS=7760000 PD=7760000
M$207 \$4 RO GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.4385e+13 AD=1.4385e+13 PS=76700000 PD=76700000
M$227 \$18 \$16 \$10 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.533e+12 AD=1.533e+12 PS=7760000 PD=7760000
M$229 \$10 DUT_Header GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.4385e+13 AD=1.4385e+13 PS=76700000 PD=76700000
M$249 \$18 RON Drain_Sense GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.533e+12 AD=1.806e+12 PS=7760000 PD=5920000
M$251 \$18 RON Drain_Force GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.806e+12 AD=1.533e+12 PS=5920000 PD=7760000
M$253 \$19 \$18 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.533e+12 AD=1.533e+12 PS=7760000 PD=7760000
M$255 \$78 GND \$23 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$256 \$79 GND \$23 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$257 \$23 \$69 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$259 \$80 GND \$69 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$260 \$81 GND \$69 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$261 \$69 \$70 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$263 \$82 GND \$70 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$264 \$83 GND \$70 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$265 \$70 \$71 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$267 \$16 RON DUT_Gate GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$268 \$84 GND \$71 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$269 \$16 RON \$17 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$270 \$85 GND \$71 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$271 \$71 \$72 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$273 \$86 GND \$72 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$274 \$87 GND \$72 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$275 \$72 \$73 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$277 \$88 GND \$73 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$278 \$89 GND \$73 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$279 \$73 \$74 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$281 \$90 GND \$74 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$282 \$91 GND \$74 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$283 \$74 \$75 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$285 \$92 GND \$75 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$286 \$93 GND \$75 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$287 \$75 \$76 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$289 \$94 GND \$76 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$290 \$95 GND \$76 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$291 \$76 OUT GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$293 \$96 GND OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$294 \$97 GND OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$295 OUT \$19 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.3335e+12 AD=1.3335e+12 PS=7570000 PD=7570000
M$297 \$19 RON GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$298 \$19 RON \$20 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
.ENDS RO_LVT_13St_x10
