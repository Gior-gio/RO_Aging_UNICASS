** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/FF/FF.sch
.subckt FF VDD D Q_N Q CLK GND
*.PININFO GND:B CLK:B VDD:B Q:B Q_N:B D:B
x1 CLKN VDD net1 D GND CLK passgate_DIV
x2 VDD net2 net1 GND inv_DIV
x3 CLK VDD net1 net4 GND CLKN passgate_DIV
x4 VDD net4 net2 GND inv_DIV
x5 CLK VDD net3 net2 GND CLKN passgate_DIV
x6 VDD net5 net3 GND inv_DIV
x7 CLKN VDD net3 Q_N GND CLK passgate_DIV
x8 VDD Q Q_N GND inv_DIV
x10 VDD CLKN CLK GND inv_DIV
x9 VDD Q_N net5 GND inv_DIV
.ends

* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/DIV/passgate_DIV/passgate_DIV.sym # of pins=6
** sym_path: /foss/designs/RO_Aging_UNICASS/DIV/passgate_DIV/passgate_DIV.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/passgate_DIV/passgate_DIV.sch
.subckt passgate_DIV CLKN VDD OUT IN GND CLK
*.PININFO VDD:B OUT:B GND:B IN:B CLKN:B CLK:B
M3 IN CLK OUT GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
M1 IN CLKN OUT VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  inv_DIV.sym # of pins=4
** sym_path: /foss/designs/RO_Aging_UNICASS/DIV/inv_DIV/inv_DIV.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/inv_DIV/inv_DIV.sch
.subckt inv_DIV VDD OUT IN GND
*.PININFO VDD:B OUT:B GND:B IN:B
M3 OUT IN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
M1 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends

.end
