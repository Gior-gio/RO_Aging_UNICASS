* Extracted by KLayout with SKY130 LVS runset on : 06/11/2024 01:14

.SUBCKT inverter VSS Out In VDD
M$1 VDD In Out VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$5 Out In VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
.ENDS inverter
