magic
tech sky130A
magscale 1 2
timestamp 1728421585
<< checkpaint >>
rect -944 -2699 1998 331
<< error_s >>
rect 129 -906 187 -900
rect 129 -940 141 -906
rect 129 -946 187 -940
rect 101 -1200 200 -1180
rect 129 -1228 187 -1208
rect 129 -1248 141 -1228
rect 129 -1254 187 -1248
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
use sky130_fd_pr__nfet_01v8_4A3DHF  XM1
timestamp 0
transform 1 0 527 0 1 -1184
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_hvt_HVTLRR  XM2
timestamp 0
transform 1 0 158 0 1 -1077
box -211 -309 211 309
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 Out
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 In
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VSS
port 3 nsew
<< end >>
