* Extracted by KLayout with SKY130 LVS runset on : 04/11/2024 04:38

.SUBCKT rovcel3_LVT GND RON RO DUT_Gate OUT IN VDD
M$1 \$74 IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$5 VDD RON \$74 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$45 OUT RO DUT_Gate VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$46 OUT RO \$16 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$47 OUT RON \$16 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$48 OUT RON DUT_Gate GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$49 GND RO \$38 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.26e+13 AD=1.26e+13 PS=96000000 PD=96000000
M$69 \$38 IN OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000 AS=1.26e+12
+ AD=1.26e+12 PS=9600000 PD=9600000
.ENDS rovcel3_LVT
