** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/rovcel4_LVT/rovcel4_LVT.sch
.subckt rovcel4_LVT VDD OUT GND RON IN
*.PININFO OUT:B RON:B IN:B GND:B VDD:B
M1 OUT IN GND GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 nf=1 m=2
M2 OUT IN net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 nf=1 m=4
M3 net1 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 nf=1 m=40
* noconn #net2
x2 VDD OUT net2 RON GND VDD passgate_LVT
x3 VDD OUT GND RON GND VDD passgate_LVT
.ends

* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/passgate_LVT/passgate_LVT.sym # of pins=6
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/passgate_LVT/passgate_LVT.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/passgate_LVT/passgate_LVT.sch
.subckt passgate_LVT CLKN IN OUT CLK GND VDD
*.PININFO CLKN:B CLK:B IN:B OUT:B VDD:B GND:B
M3 IN CLK OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 nf=1 m=1
M1 IN CLKN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 nf=1 m=1
.ends

.end
