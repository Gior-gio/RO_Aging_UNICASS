magic
tech sky130
timestamp 1729529908
<< checkpaint >>
<< l67d20 >>
<< l68d20 >>
<< l67d44 >>
<< end >>
