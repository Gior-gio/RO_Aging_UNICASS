** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/rovcel2_LVT/rovcel2_LVT.sch
.subckt rovcel2_LVT VDD GND IN OUT
*.PININFO OUT:B IN:B VDD:B GND:B
* noconn #net1
* noconn #net2
x1 VDD IN OUT GND inv_LVT
x2 VDD OUT net1 GND GND VDD passgate_LVT
x3 VDD OUT net2 GND GND VDD passgate_LVT
.ends

* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/inv_LVT/inv_LVT.sym # of pins=4
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/inv_LVT/inv_LVT.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/inv_LVT/inv_LVT.sch
.subckt inv_LVT VDD IN OUT GND
*.PININFO VDD:B IN:B OUT:B GND:B
M1 OUT IN GND GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 nf=1 m=2
M2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 nf=1 m=4
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/passgate_LVT/passgate_LVT.sym # of pins=6
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/passgate_LVT/passgate_LVT.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/passgate_LVT/passgate_LVT.sch
.subckt passgate_LVT CLKN IN OUT CLK GND VDD
*.PININFO CLKN:B CLK:B IN:B OUT:B VDD:B GND:B
M3 IN CLK OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 nf=1 m=1
M1 IN CLKN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 nf=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
