magic
tech sky130A
timestamp 1727311909
<< properties >>
string (UNNAMED) gencell
<< end >>
