* Extracted by KLayout with SKY130 LVS runset on : 05/11/2024 01:55

.SUBCKT rovcel1_x1_LVT GND DUT_Footer DUT_Header Drain_Sense Drain\x20Force IN
+ VDD
M$1 \$81 IN \$8 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$5 VDD DUT_Footer \$81 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$45 \$8 \$15 Drain_Sense VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$49 \$8 \$15 Drain\x20Force VDD sky130_fd_pr__pfet_01v8_lvt L=350000
+ W=19000000 AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$53 GND DUT_Header \$9 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.26e+13 AD=1.26e+13 PS=96000000 PD=96000000
M$73 \$8 \$20 Drain_Sense GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$74 Drain\x20Force \$20 \$8 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$75 \$9 IN \$8 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000 AS=1.26e+12
+ AD=1.26e+12 PS=9600000 PD=9600000
.ENDS rovcel1_x1_LVT
