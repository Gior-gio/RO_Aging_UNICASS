magic
tech sky130
timestamp 1729529908
<< checkpaint >>
rect 1 -1 3 3
<< l68d20 >>
<< l66d44 >>
rect 1 -1 2 0
rect 1 2 2 3
<< l69d20 >>
<< l68d16 >>
rect 1 2 2 3
rect 1 -1 2 0
<< l69d16 >>
<< labels >>
rlabel l68d5 1.56 2.275 1.56 2.275 0 VDD
rlabel l68d5 1.88 0.95 1.88 0.95 0 In
rlabel l68d5 1.56 -0.355 1.56 -0.355 0 VSS
rlabel l69d5 2.215 0.925 2.215 0.925 0 Out
use pfet pfet_1
timestamp 1729529908
transform -1 0 2 0 1 2
box 0 -1 1 1
use vias_genx241 vias_genx241_1
timestamp 1729529908
transform 1 0 2 0 1 -1
box 0 0 0 1
use vias_genx241 vias_genx241_2
timestamp 1729529908
transform 1 0 2 0 1 2
box 0 0 0 1
use vias_genx242 vias_genx242_1
timestamp 1729529908
transform 1 0 1 0 1 -1
box 0 0 0 1
use vias_genx242 vias_genx242_2
timestamp 1729529908
transform 1 0 1 0 1 2
box 0 0 0 1
use nfet nfet_1
timestamp 1729529908
transform -1 0 2 0 1 -1
box 0 0 1 2
<< end >>
