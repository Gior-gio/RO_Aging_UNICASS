* Extracted by KLayout with SKY130 LVS runset on : 04/11/2024 05:27

.SUBCKT rovcel4_LVT GND RON OUT IN VDD
M$1 \$28 IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$5 VDD RON \$28 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$45 OUT VDD GND VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$46 OUT VDD \$11 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$47 OUT RON \$11 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$48 OUT RON GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$49 GND IN OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000 AS=1.26e+12
+ AD=1.26e+12 PS=9600000 PD=9600000
.ENDS rovcel4_LVT
