* Extracted by KLayout with SKY130 LVS runset on : 09/11/2024 21:29

.SUBCKT FF CLK GND Q_N Q D VDD
M$1 VDD Q_N Q VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000 AS=600000000000
+ AD=600000000000 PS=5200000 PD=5200000
M$2 \$6 CLK \$13 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$3 Q_N \$15 VDD VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000 AS=600000000000
+ AD=600000000000 PS=5200000 PD=5200000
M$4 VDD \$14 \$15 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$7 Q_N \$1 \$14 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$9 VDD CLK \$1 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000 AS=600000000000
+ AD=600000000000 PS=5200000 PD=5200000
M$10 \$5 \$13 VDD VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$11 \$5 CLK \$14 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$12 D \$1 \$13 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$15 VDD \$5 \$6 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000 AS=600000000000
+ AD=600000000000 PS=5200000 PD=5200000
M$17 GND \$13 \$5 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$18 GND CLK \$1 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$19 Q_N CLK \$14 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000 AS=195000000000
+ AD=195000000000 PS=1900000 PD=1900000
M$20 GND Q_N Q GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$21 D CLK \$13 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000 AS=195000000000
+ AD=195000000000 PS=1900000 PD=1900000
M$22 GND \$15 Q_N GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$23 \$6 \$1 \$13 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000 AS=195000000000
+ AD=195000000000 PS=1900000 PD=1900000
M$24 GND \$14 \$15 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$25 GND \$5 \$6 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$26 \$5 \$1 \$14 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000 AS=195000000000
+ AD=195000000000 PS=1900000 PD=1900000
.ENDS FF
