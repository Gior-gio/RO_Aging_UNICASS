magic
tech sky130
timestamp 1729529908
<< checkpaint >>
rect 0 0 1 2
<< l67d20 >>
<< l68d20 >>
rect 0 0 1 1
<< l67d44 >>
<< l65d20 >>
rect 0 0 1 1
<< l66d44 >>
<< l66d20 >>
rect 0 1 1 2
<< l95d20 >>
rect 0 1 1 2
<< l65d44 >>
<< l94d20 >>
<< l93d44 >>
rect 0 0 1 1
<< end >>
