* Extracted by KLayout with SKY130 LVS runset on : 06/11/2024 05:40

.SUBCKT RingOscilator_hvt_13_x10 DRAIN_SENSE DRAIN_FORCE DUT_FOOTER DUT_GATE
+ DUT_HEADER NOT_RO_CON RO_CON VSS VDD A[1]
X$8 VSS DUT_HEADER \$42 \$37 VDD DUT_FOOTER rovcel
X$10 NOT_RO_CON \$37 DUT_GATE RO_CON VDD VSS passGate_hvt
X$13 VSS RO_CON \$37 \$20 VDD NOT_RO_CON rovcel
X$23 NOT_RO_CON \$37 \$I64 RO_CON VDD VSS passGate_hvt
X$25 NOT_RO_CON \$27 \$I66 VDD VDD VSS passGate_hvt
X$27 NOT_RO_CON \$27 VSS VDD VDD VSS passGate_hvt
M$1 VDD NOT_RO_CON \$I98 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=190000000
+ AS=6.25575e+13 AD=6.25575e+13 PS=221090000 PD=221090000
M$41 \$I98 \$42 \$27 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$45 \$27 \$42 VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
M$47 \$42 RO_CON DRAIN_SENSE VDD sky130_fd_pr__pfet_01v8_hvt L=150000
+ W=19000000 AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$51 DRAIN_SENSE NOT_RO_CON \$42 VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000
+ AS=1.323e+12 AD=1.323e+12 PS=7560000 PD=7560000
M$53 \$42 RO_CON DRAIN_FORCE VDD sky130_fd_pr__pfet_01v8_hvt L=150000
+ W=190000000 AS=6.4588125e+13 AD=6.5181875e+13 PS=221945000 PD=222195000
M$93 DRAIN_FORCE NOT_RO_CON \$42 VSS sky130_fd_pr__nfet_01v8 L=150000
+ W=42000000 AS=1.3797e+13 AD=1.3797e+13 PS=57240000 PD=57240000
M$113 VDD A[1] \$I19 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$117 \$I19 A[1] VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000
+ AS=1.323e+12 AD=1.323e+12 PS=7560000 PD=7560000
M$119 VDD \$27 A[1] VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$123 A[1] \$27 VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
M$125 VDD \$I19 \$I10 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$129 \$I10 \$I19 VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000
+ AS=1.323e+12 AD=1.323e+12 PS=7560000 PD=7560000
M$131 VDD \$I10 \$I17 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$135 \$I17 \$I10 VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000
+ AS=1.323e+12 AD=1.323e+12 PS=7560000 PD=7560000
M$137 VDD \$I17 \$I15 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$141 \$I15 \$I17 VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000
+ AS=1.323e+12 AD=1.323e+12 PS=7560000 PD=7560000
M$143 VDD \$I15 \$I18 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$147 \$I18 \$I15 VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000
+ AS=1.323e+12 AD=1.323e+12 PS=7560000 PD=7560000
M$149 VDD \$I18 \$I14 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$153 \$I14 \$I18 VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000
+ AS=1.323e+12 AD=1.323e+12 PS=7560000 PD=7560000
M$155 VDD \$I14 \$I13 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$159 \$I13 \$I14 VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000
+ AS=1.323e+12 AD=1.323e+12 PS=7560000 PD=7560000
M$161 VDD \$I13 \$I12 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$165 \$I12 \$I13 VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000
+ AS=1.323e+12 AD=1.323e+12 PS=7560000 PD=7560000
M$167 VDD \$I12 \$20 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$171 \$20 \$I12 VSS VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000
+ AS=1.323e+12 AD=1.323e+12 PS=7560000 PD=7560000
M$173 \$I19 VDD \$I107 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$174 \$I19 VDD \$I106 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$175 A[1] VDD \$I111 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$176 A[1] VDD \$I110 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$177 \$I10 VDD \$I115 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$178 \$I10 VDD \$I114 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$179 \$I17 VDD \$I119 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$180 \$I17 VDD \$I118 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$181 \$I15 VDD \$I123 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$182 \$I15 VDD \$I122 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$183 \$I18 VDD \$I127 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$184 \$I18 VDD \$I126 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$185 \$I14 VDD \$I131 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$186 \$I14 VDD \$I130 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$187 \$I13 VDD \$I135 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$188 \$I13 VDD \$I134 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$189 \$I12 VDD \$I139 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$190 \$I12 VDD \$I138 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$191 \$20 VDD \$I143 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$192 \$20 VDD \$I142 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$193 \$I19 VSS \$I107 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$194 \$I19 VSS \$I106 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$195 A[1] VSS \$I111 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$196 A[1] VSS \$I110 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$197 \$I10 VSS \$I115 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$198 \$I10 VSS \$I114 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$199 \$I17 VSS \$I119 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$200 \$I17 VSS \$I118 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$201 \$I15 VSS \$I123 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$202 \$I15 VSS \$I122 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$203 \$I18 VSS \$I127 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$204 \$I18 VSS \$I126 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$205 \$I14 VSS \$I131 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$206 \$I14 VSS \$I130 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$207 \$I13 VSS \$I135 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$208 \$I13 VSS \$I134 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$209 \$I12 VSS \$I139 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$210 \$I12 VSS \$I138 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$211 \$20 VSS \$I143 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$212 \$20 VSS \$I142 VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
.ENDS RingOscilator_hvt_13_x10

.SUBCKT passGate_hvt CLK In Out CLKN VDD VSS
M$1 In CLKN Out VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$2 In CLK Out VSS sky130_fd_pr__nfet_01v8 L=150000 W=450000 AS=135000000000
+ AD=135000000000 PS=1500000 PD=1500000
.ENDS passGate_hvt

.SUBCKT rovcel VSS N Out IN VDD P
M$1 VDD P \$79 VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=190000000
+ AS=6.25575e+13 AD=6.25575e+13 PS=221090000 PD=221090000
M$41 \$79 IN Out VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=19000000
+ AS=6.1275e+12 AD=6.1275e+12 PS=26330000 PD=26330000
M$45 VSS N \$9 VSS sky130_fd_pr__nfet_01v8 L=150000 W=42000000 AS=1.3797e+13
+ AD=1.3797e+13 PS=57240000 PD=57240000
M$65 Out IN \$9 VSS sky130_fd_pr__nfet_01v8 L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
.ENDS rovcel
