magic
tech sky130A
magscale 1 2
timestamp 1728409320
<< error_p >>
rect -29 126 29 132
rect -29 92 -17 126
rect -29 86 29 92
rect -29 -92 29 -86
rect -29 -126 -17 -92
rect -29 -132 29 -126
<< nwell >>
rect -211 -264 211 264
<< pmoshvt >>
rect -15 -45 15 45
<< pdiff >>
rect -73 33 -15 45
rect -73 -33 -61 33
rect -27 -33 -15 33
rect -73 -45 -15 -33
rect 15 33 73 45
rect 15 -33 27 33
rect 61 -33 73 33
rect 15 -45 73 -33
<< pdiffc >>
rect -61 -33 -27 33
rect 27 -33 61 33
<< nsubdiff >>
rect -175 194 -79 228
rect 79 194 175 228
rect -175 132 -141 194
rect 141 132 175 194
rect -175 -194 -141 -132
rect 141 -194 175 -132
rect -175 -228 -79 -194
rect 79 -228 175 -194
<< nsubdiffcont >>
rect -79 194 79 228
rect -175 -132 -141 132
rect 141 -132 175 132
rect -79 -228 79 -194
<< poly >>
rect -33 126 33 142
rect -33 92 -17 126
rect 17 92 33 126
rect -33 76 33 92
rect -15 45 15 76
rect -15 -76 15 -45
rect -33 -92 33 -76
rect -33 -126 -17 -92
rect 17 -126 33 -92
rect -33 -142 33 -126
<< polycont >>
rect -17 92 17 126
rect -17 -126 17 -92
<< locali >>
rect -175 194 -79 228
rect 79 194 175 228
rect -175 132 -141 194
rect 141 132 175 194
rect -33 92 -17 126
rect 17 92 33 126
rect -61 33 -27 49
rect -61 -49 -27 -33
rect 27 33 61 49
rect 27 -49 61 -33
rect -33 -126 -17 -92
rect 17 -126 33 -92
rect -175 -194 -141 -132
rect 141 -194 175 -132
rect -175 -228 -79 -194
rect 79 -228 175 -194
<< viali >>
rect -17 92 17 126
rect -61 -33 -27 33
rect 27 -33 61 33
rect -17 -126 17 -92
<< metal1 >>
rect -29 126 29 132
rect -29 92 -17 126
rect 17 92 29 126
rect -29 86 29 92
rect -67 33 -21 45
rect -67 -33 -61 33
rect -27 -33 -21 33
rect -67 -45 -21 -33
rect 21 33 67 45
rect 21 -33 27 33
rect 61 -33 67 33
rect 21 -45 67 -33
rect -29 -92 29 -86
rect -29 -126 -17 -92
rect 17 -126 29 -92
rect -29 -132 29 -126
<< properties >>
string FIXED_BBOX -158 -211 158 211
string gencell sky130_fd_pr__pfet_01v8_hvt
string library sky130
string parameters w 0.45 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 1
<< end >>
