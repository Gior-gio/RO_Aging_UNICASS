* Extracted by KLayout with SKY130 LVS runset on : 03/11/2024 02:05

.SUBCKT rovcel VSS N Out IN VDD P
M$1 VDD P \$72 VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=190 AS=62.5575
+ AD=62.5575 PS=221.09 PD=221.09
M$41 \$72 IN Out VDD sky130_fd_pr__pfet_01v8_hvt L=0.15 W=19 AS=6.1275
+ AD=6.1275 PS=26.33 PD=26.33
M$45 VSS N \$6 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=37.8 AS=12.411 AD=12.411
+ PS=51.72 PD=51.72
M$63 Out IN \$6 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=4.2 AS=1.323 AD=1.323
+ PS=7.56 PD=7.56
.ENDS rovcel
