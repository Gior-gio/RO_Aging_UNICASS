* Extracted by KLayout with SKY130 LVS runset on : 03/11/2024 20:20

.SUBCKT nmos_lvt VG VD VSS
M$1 VD VG \$3 VSS sky130_fd_pr__nfet_01v8_lvt L=150000 W=4200000 AS=1.323e+12
+ AD=1.323e+12 PS=7560000 PD=7560000
.ENDS nmos_lvt
