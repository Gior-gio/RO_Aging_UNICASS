* Extracted by KLayout with SKY130 LVS runset on : 03/11/2024 23:28

.SUBCKT passGate_lvt CLKN CLK OUT IN VDD GND
M$1 IN CLK OUT GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$2 IN CLKN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
.ENDS passGate_lvt
