* Extracted by KLayout with SKY130 LVS runset on : 05/11/2024 14:50

.SUBCKT load_x10 VSS Out In A VDD AB
M$1 In AB Out VDD sky130_fd_pr__pfet_01v8_hvt L=150000 W=190000000
+ AS=6.4588125e+13 AD=6.5181875e+13 PS=221945000 PD=222195000
M$41 Out A In VSS sky130_fd_pr__nfet_01v8 L=150000 W=42000000 AS=1.3797e+13
+ AD=1.3797e+13 PS=57240000 PD=57240000
.ENDS load_x10
