* Extracted by KLayout with SKY130 LVS runset on : 05/11/2024 15:34

.SUBCKT vias_gen$10$2$1$1$1$1$1$1
.ENDS vias_gen$10$2$1$1$1$1$1$1

.SUBCKT vias_gen$2$1$2$1$1$1$1$1$1
.ENDS vias_gen$2$1$2$1$1$1$1$1$1

.SUBCKT pfet$2$2$1$1$1$1$1$1
.ENDS pfet$2$2$1$1$1$1$1$1

.SUBCKT vias_gen$6$2$1$1$1$1$1$1
.ENDS vias_gen$6$2$1$1$1$1$1$1

.SUBCKT vias_gen$18$2$1$1$1$1$1$1
.ENDS vias_gen$18$2$1$1$1$1$1$1

.SUBCKT nfet$2$2$1$1$1$1$1$1
.ENDS nfet$2$2$1$1$1$1$1$1

.SUBCKT vias_gen$7$2$1$1$1$1$1$1
.ENDS vias_gen$7$2$1$1$1$1$1$1

.SUBCKT vias_gen$10$1$1$1$1$1$1$1$1
.ENDS vias_gen$10$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$2$1$1$1$1$1$1$1$1$1
.ENDS vias_gen$2$1$1$1$1$1$1$1$1$1

.SUBCKT pfet$2$1$1$1$1$1$1$1$1
.ENDS pfet$2$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$6$1$1$1$1$1$1$1$1
.ENDS vias_gen$6$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$18$1$1$1$1$1$1$1$1
.ENDS vias_gen$18$1$1$1$1$1$1$1$1

.SUBCKT nfet$2$1$1$1$1$1$1$1$1
.ENDS nfet$2$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$7$1$1$1$1$1$1$1$1
.ENDS vias_gen$7$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$10$3$1$1$1$1$1
.ENDS vias_gen$10$3$1$1$1$1$1

.SUBCKT vias_gen$2$1$3$1$1$1$1$1
.ENDS vias_gen$2$1$3$1$1$1$1$1

.SUBCKT pfet$2$3$1$1$1$1$1
.ENDS pfet$2$3$1$1$1$1$1

.SUBCKT vias_gen$6$3$1$1$1$1$1
.ENDS vias_gen$6$3$1$1$1$1$1

.SUBCKT vias_gen$18$3$1$1$1$1$1
.ENDS vias_gen$18$3$1$1$1$1$1

.SUBCKT nfet$2$3$1$1$1$1$1
.ENDS nfet$2$3$1$1$1$1$1

.SUBCKT vias_gen$7$3$1$1$1$1$1
.ENDS vias_gen$7$3$1$1$1$1$1

.SUBCKT vias_gen$10$1$2$1$1$1$1$1
.ENDS vias_gen$10$1$2$1$1$1$1$1

.SUBCKT vias_gen$2$1$1$2$1$1$1$1$1
.ENDS vias_gen$2$1$1$2$1$1$1$1$1

.SUBCKT pfet$2$1$2$1$1$1$1$1
.ENDS pfet$2$1$2$1$1$1$1$1

.SUBCKT vias_gen$6$1$2$1$1$1$1$1
.ENDS vias_gen$6$1$2$1$1$1$1$1

.SUBCKT vias_gen$18$1$2$1$1$1$1$1
.ENDS vias_gen$18$1$2$1$1$1$1$1

.SUBCKT nfet$2$1$2$1$1$1$1$1
.ENDS nfet$2$1$2$1$1$1$1$1

.SUBCKT vias_gen$7$1$2$1$1$1$1$1
.ENDS vias_gen$7$1$2$1$1$1$1$1

.SUBCKT vias_gen$10$2$2$1$1$1$1
.ENDS vias_gen$10$2$2$1$1$1$1

.SUBCKT vias_gen$2$1$2$2$1$1$1$1
.ENDS vias_gen$2$1$2$2$1$1$1$1

.SUBCKT pfet$2$2$2$1$1$1$1
.ENDS pfet$2$2$2$1$1$1$1

.SUBCKT vias_gen$6$2$2$1$1$1$1
.ENDS vias_gen$6$2$2$1$1$1$1

.SUBCKT vias_gen$18$2$2$1$1$1$1
.ENDS vias_gen$18$2$2$1$1$1$1

.SUBCKT nfet$2$2$2$1$1$1$1
.ENDS nfet$2$2$2$1$1$1$1

.SUBCKT vias_gen$7$2$2$1$1$1$1
.ENDS vias_gen$7$2$2$1$1$1$1

.SUBCKT vias_gen$10$1$1$2$1$1$1$1
.ENDS vias_gen$10$1$1$2$1$1$1$1

.SUBCKT vias_gen$2$1$1$1$2$1$1$1$1
.ENDS vias_gen$2$1$1$1$2$1$1$1$1

.SUBCKT pfet$2$1$1$2$1$1$1$1
.ENDS pfet$2$1$1$2$1$1$1$1

.SUBCKT vias_gen$6$1$1$2$1$1$1$1
.ENDS vias_gen$6$1$1$2$1$1$1$1

.SUBCKT vias_gen$18$1$1$2$1$1$1$1
.ENDS vias_gen$18$1$1$2$1$1$1$1

.SUBCKT nfet$2$1$1$2$1$1$1$1
.ENDS nfet$2$1$1$2$1$1$1$1

.SUBCKT vias_gen$7$1$1$2$1$1$1$1
.ENDS vias_gen$7$1$1$2$1$1$1$1

.SUBCKT vias_gen$10$2$1$2$1$1$1
.ENDS vias_gen$10$2$1$2$1$1$1

.SUBCKT vias_gen$2$1$2$1$2$1$1$1
.ENDS vias_gen$2$1$2$1$2$1$1$1

.SUBCKT pfet$2$2$1$2$1$1$1
.ENDS pfet$2$2$1$2$1$1$1

.SUBCKT vias_gen$6$2$1$2$1$1$1
.ENDS vias_gen$6$2$1$2$1$1$1

.SUBCKT vias_gen$18$2$1$2$1$1$1
.ENDS vias_gen$18$2$1$2$1$1$1

.SUBCKT nfet$2$2$1$2$1$1$1
.ENDS nfet$2$2$1$2$1$1$1

.SUBCKT vias_gen$7$2$1$2$1$1$1
.ENDS vias_gen$7$2$1$2$1$1$1

.SUBCKT vias_gen$10$1$1$1$2$1$1$1
.ENDS vias_gen$10$1$1$1$2$1$1$1

.SUBCKT vias_gen$2$1$1$1$1$2$1$1$1
.ENDS vias_gen$2$1$1$1$1$2$1$1$1

.SUBCKT pfet$2$1$1$1$2$1$1$1
.ENDS pfet$2$1$1$1$2$1$1$1

.SUBCKT vias_gen$6$1$1$1$2$1$1$1
.ENDS vias_gen$6$1$1$1$2$1$1$1

.SUBCKT vias_gen$18$1$1$1$2$1$1$1
.ENDS vias_gen$18$1$1$1$2$1$1$1

.SUBCKT nfet$2$1$1$1$2$1$1$1
.ENDS nfet$2$1$1$1$2$1$1$1

.SUBCKT vias_gen$7$1$1$1$2$1$1$1
.ENDS vias_gen$7$1$1$1$2$1$1$1

.SUBCKT vias_gen$10$3$2$1$1$1
.ENDS vias_gen$10$3$2$1$1$1

.SUBCKT vias_gen$2$1$3$2$1$1$1
.ENDS vias_gen$2$1$3$2$1$1$1

.SUBCKT pfet$2$3$2$1$1$1
.ENDS pfet$2$3$2$1$1$1

.SUBCKT vias_gen$6$3$2$1$1$1
.ENDS vias_gen$6$3$2$1$1$1

.SUBCKT vias_gen$18$3$2$1$1$1
.ENDS vias_gen$18$3$2$1$1$1

.SUBCKT nfet$2$3$2$1$1$1
.ENDS nfet$2$3$2$1$1$1

.SUBCKT vias_gen$7$3$2$1$1$1
.ENDS vias_gen$7$3$2$1$1$1

.SUBCKT vias_gen$10$1$2$2$1$1$1
.ENDS vias_gen$10$1$2$2$1$1$1

.SUBCKT vias_gen$2$1$1$2$2$1$1$1
.ENDS vias_gen$2$1$1$2$2$1$1$1

.SUBCKT pfet$2$1$2$2$1$1$1
.ENDS pfet$2$1$2$2$1$1$1

.SUBCKT vias_gen$6$1$2$2$1$1$1
.ENDS vias_gen$6$1$2$2$1$1$1

.SUBCKT vias_gen$18$1$2$2$1$1$1
.ENDS vias_gen$18$1$2$2$1$1$1

.SUBCKT nfet$2$1$2$2$1$1$1
.ENDS nfet$2$1$2$2$1$1$1

.SUBCKT vias_gen$7$1$2$2$1$1$1
.ENDS vias_gen$7$1$2$2$1$1$1

.SUBCKT vias_gen$10$2$1$1$1$2$1
.ENDS vias_gen$10$2$1$1$1$2$1

.SUBCKT vias_gen$2$1$2$1$1$1$2$1
.ENDS vias_gen$2$1$2$1$1$1$2$1

.SUBCKT pfet$2$2$1$1$1$2$1
.ENDS pfet$2$2$1$1$1$2$1

.SUBCKT vias_gen$6$2$1$1$1$2$1
.ENDS vias_gen$6$2$1$1$1$2$1

.SUBCKT vias_gen$18$2$1$1$1$2$1
.ENDS vias_gen$18$2$1$1$1$2$1

.SUBCKT nfet$2$2$1$1$1$2$1
.ENDS nfet$2$2$1$1$1$2$1

.SUBCKT vias_gen$7$2$1$1$1$2$1
.ENDS vias_gen$7$2$1$1$1$2$1

.SUBCKT vias_gen$10$1$1$1$1$1$2$1
.ENDS vias_gen$10$1$1$1$1$1$2$1

.SUBCKT vias_gen$2$1$1$1$1$1$1$2$1
.ENDS vias_gen$2$1$1$1$1$1$1$2$1

.SUBCKT pfet$2$1$1$1$1$1$2$1
.ENDS pfet$2$1$1$1$1$1$2$1

.SUBCKT vias_gen$6$1$1$1$1$1$2$1
.ENDS vias_gen$6$1$1$1$1$1$2$1

.SUBCKT vias_gen$18$1$1$1$1$1$2$1
.ENDS vias_gen$18$1$1$1$1$1$2$1

.SUBCKT nfet$2$1$1$1$1$1$2$1
.ENDS nfet$2$1$1$1$1$1$2$1

.SUBCKT vias_gen$7$1$1$1$1$1$2$1
.ENDS vias_gen$7$1$1$1$1$1$2$1

.SUBCKT vias_gen$10$3$1$1$2$1
.ENDS vias_gen$10$3$1$1$2$1

.SUBCKT vias_gen$2$1$3$1$1$2$1
.ENDS vias_gen$2$1$3$1$1$2$1

.SUBCKT pfet$2$3$1$1$2$1
.ENDS pfet$2$3$1$1$2$1

.SUBCKT vias_gen$6$3$1$1$2$1
.ENDS vias_gen$6$3$1$1$2$1

.SUBCKT vias_gen$18$3$1$1$2$1
.ENDS vias_gen$18$3$1$1$2$1

.SUBCKT nfet$2$3$1$1$2$1
.ENDS nfet$2$3$1$1$2$1

.SUBCKT vias_gen$7$3$1$1$2$1
.ENDS vias_gen$7$3$1$1$2$1

.SUBCKT vias_gen$10$1$2$1$1$2$1
.ENDS vias_gen$10$1$2$1$1$2$1

.SUBCKT vias_gen$2$1$1$2$1$1$2$1
.ENDS vias_gen$2$1$1$2$1$1$2$1

.SUBCKT pfet$2$1$2$1$1$2$1
.ENDS pfet$2$1$2$1$1$2$1

.SUBCKT vias_gen$6$1$2$1$1$2$1
.ENDS vias_gen$6$1$2$1$1$2$1

.SUBCKT vias_gen$18$1$2$1$1$2$1
.ENDS vias_gen$18$1$2$1$1$2$1

.SUBCKT nfet$2$1$2$1$1$2$1
.ENDS nfet$2$1$2$1$1$2$1

.SUBCKT vias_gen$7$1$2$1$1$2$1
.ENDS vias_gen$7$1$2$1$1$2$1

.SUBCKT vias_gen$10$2$2$1$2$1
.ENDS vias_gen$10$2$2$1$2$1

.SUBCKT vias_gen$2$1$2$2$1$2$1
.ENDS vias_gen$2$1$2$2$1$2$1

.SUBCKT pfet$2$2$2$1$2$1
.ENDS pfet$2$2$2$1$2$1

.SUBCKT vias_gen$6$2$2$1$2$1
.ENDS vias_gen$6$2$2$1$2$1

.SUBCKT vias_gen$18$2$2$1$2$1
.ENDS vias_gen$18$2$2$1$2$1

.SUBCKT nfet$2$2$2$1$2$1
.ENDS nfet$2$2$2$1$2$1

.SUBCKT vias_gen$7$2$2$1$2$1
.ENDS vias_gen$7$2$2$1$2$1

.SUBCKT vias_gen$10$1$1$2$1$2$1
.ENDS vias_gen$10$1$1$2$1$2$1

.SUBCKT vias_gen$2$1$1$1$2$1$2$1
.ENDS vias_gen$2$1$1$1$2$1$2$1

.SUBCKT pfet$2$1$1$2$1$2$1
.ENDS pfet$2$1$1$2$1$2$1

.SUBCKT vias_gen$6$1$1$2$1$2$1
.ENDS vias_gen$6$1$1$2$1$2$1

.SUBCKT vias_gen$18$1$1$2$1$2$1
.ENDS vias_gen$18$1$1$2$1$2$1

.SUBCKT nfet$2$1$1$2$1$2$1
.ENDS nfet$2$1$1$2$1$2$1

.SUBCKT vias_gen$7$1$1$2$1$2$1
.ENDS vias_gen$7$1$1$2$1$2$1

.SUBCKT vias_gen$10$2$1$2$2$1
.ENDS vias_gen$10$2$1$2$2$1

.SUBCKT vias_gen$2$1$2$1$2$2$1
.ENDS vias_gen$2$1$2$1$2$2$1

.SUBCKT pfet$2$2$1$2$2$1
.ENDS pfet$2$2$1$2$2$1

.SUBCKT vias_gen$6$2$1$2$2$1
.ENDS vias_gen$6$2$1$2$2$1

.SUBCKT vias_gen$18$2$1$2$2$1
.ENDS vias_gen$18$2$1$2$2$1

.SUBCKT nfet$2$2$1$2$2$1
.ENDS nfet$2$2$1$2$2$1

.SUBCKT vias_gen$7$2$1$2$2$1
.ENDS vias_gen$7$2$1$2$2$1

.SUBCKT vias_gen$10$1$1$1$2$2$1
.ENDS vias_gen$10$1$1$1$2$2$1

.SUBCKT vias_gen$2$1$1$1$1$2$2$1
.ENDS vias_gen$2$1$1$1$1$2$2$1

.SUBCKT pfet$2$1$1$1$2$2$1
.ENDS pfet$2$1$1$1$2$2$1

.SUBCKT vias_gen$6$1$1$1$2$2$1
.ENDS vias_gen$6$1$1$1$2$2$1

.SUBCKT vias_gen$18$1$1$1$2$2$1
.ENDS vias_gen$18$1$1$1$2$2$1

.SUBCKT nfet$2$1$1$1$2$2$1
.ENDS nfet$2$1$1$1$2$2$1

.SUBCKT vias_gen$7$1$1$1$2$2$1
.ENDS vias_gen$7$1$1$1$2$2$1

.SUBCKT vias_gen$10$3$2$2$1
.ENDS vias_gen$10$3$2$2$1

.SUBCKT vias_gen$2$1$3$2$2$1
.ENDS vias_gen$2$1$3$2$2$1

.SUBCKT pfet$2$3$2$2$1
.ENDS pfet$2$3$2$2$1

.SUBCKT vias_gen$6$3$2$2$1
.ENDS vias_gen$6$3$2$2$1

.SUBCKT vias_gen$18$3$2$2$1
.ENDS vias_gen$18$3$2$2$1

.SUBCKT nfet$2$3$2$2$1
.ENDS nfet$2$3$2$2$1

.SUBCKT vias_gen$7$3$2$2$1
.ENDS vias_gen$7$3$2$2$1

.SUBCKT vias_gen$10$1$2$2$2$1
.ENDS vias_gen$10$1$2$2$2$1

.SUBCKT vias_gen$2$1$1$2$2$2$1
.ENDS vias_gen$2$1$1$2$2$2$1

.SUBCKT pfet$2$1$2$2$2$1
.ENDS pfet$2$1$2$2$2$1

.SUBCKT vias_gen$6$1$2$2$2$1
.ENDS vias_gen$6$1$2$2$2$1

.SUBCKT vias_gen$18$1$2$2$2$1
.ENDS vias_gen$18$1$2$2$2$1

.SUBCKT nfet$2$1$2$2$2$1
.ENDS nfet$2$1$2$2$2$1

.SUBCKT vias_gen$7$1$2$2$2$1
.ENDS vias_gen$7$1$2$2$2$1

.SUBCKT vias_gen$10$2$1$1$1$1$2
.ENDS vias_gen$10$2$1$1$1$1$2

.SUBCKT vias_gen$2$1$2$1$1$1$1$2
.ENDS vias_gen$2$1$2$1$1$1$1$2

.SUBCKT pfet$2$2$1$1$1$1$2
.ENDS pfet$2$2$1$1$1$1$2

.SUBCKT vias_gen$6$2$1$1$1$1$2
.ENDS vias_gen$6$2$1$1$1$1$2

.SUBCKT vias_gen$18$2$1$1$1$1$2
.ENDS vias_gen$18$2$1$1$1$1$2

.SUBCKT nfet$2$2$1$1$1$1$2
.ENDS nfet$2$2$1$1$1$1$2

.SUBCKT vias_gen$7$2$1$1$1$1$2
.ENDS vias_gen$7$2$1$1$1$1$2

.SUBCKT vias_gen$10$1$1$1$1$1$1$2
.ENDS vias_gen$10$1$1$1$1$1$1$2

.SUBCKT vias_gen$2$1$1$1$1$1$1$1$2
.ENDS vias_gen$2$1$1$1$1$1$1$1$2

.SUBCKT pfet$2$1$1$1$1$1$1$2
.ENDS pfet$2$1$1$1$1$1$1$2

.SUBCKT vias_gen$6$1$1$1$1$1$1$2
.ENDS vias_gen$6$1$1$1$1$1$1$2

.SUBCKT vias_gen$18$1$1$1$1$1$1$2
.ENDS vias_gen$18$1$1$1$1$1$1$2

.SUBCKT nfet$2$1$1$1$1$1$1$2
.ENDS nfet$2$1$1$1$1$1$1$2

.SUBCKT vias_gen$7$1$1$1$1$1$1$2
.ENDS vias_gen$7$1$1$1$1$1$1$2

.SUBCKT vias_gen$10$3$1$1$1$2
.ENDS vias_gen$10$3$1$1$1$2

.SUBCKT vias_gen$2$1$3$1$1$1$2
.ENDS vias_gen$2$1$3$1$1$1$2

.SUBCKT pfet$2$3$1$1$1$2
.ENDS pfet$2$3$1$1$1$2

.SUBCKT vias_gen$6$3$1$1$1$2
.ENDS vias_gen$6$3$1$1$1$2

.SUBCKT vias_gen$18$3$1$1$1$2
.ENDS vias_gen$18$3$1$1$1$2

.SUBCKT nfet$2$3$1$1$1$2
.ENDS nfet$2$3$1$1$1$2

.SUBCKT vias_gen$7$3$1$1$1$2
.ENDS vias_gen$7$3$1$1$1$2

.SUBCKT vias_gen$10$1$2$1$1$1$2
.ENDS vias_gen$10$1$2$1$1$1$2

.SUBCKT vias_gen$2$1$1$2$1$1$1$2
.ENDS vias_gen$2$1$1$2$1$1$1$2

.SUBCKT pfet$2$1$2$1$1$1$2
.ENDS pfet$2$1$2$1$1$1$2

.SUBCKT vias_gen$6$1$2$1$1$1$2
.ENDS vias_gen$6$1$2$1$1$1$2

.SUBCKT vias_gen$18$1$2$1$1$1$2
.ENDS vias_gen$18$1$2$1$1$1$2

.SUBCKT nfet$2$1$2$1$1$1$2
.ENDS nfet$2$1$2$1$1$1$2

.SUBCKT vias_gen$7$1$2$1$1$1$2
.ENDS vias_gen$7$1$2$1$1$1$2

.SUBCKT vias_gen$10$2$2$1$1$2
.ENDS vias_gen$10$2$2$1$1$2

.SUBCKT vias_gen$2$1$2$2$1$1$2
.ENDS vias_gen$2$1$2$2$1$1$2

.SUBCKT pfet$2$2$2$1$1$2
.ENDS pfet$2$2$2$1$1$2

.SUBCKT vias_gen$6$2$2$1$1$2
.ENDS vias_gen$6$2$2$1$1$2

.SUBCKT vias_gen$18$2$2$1$1$2
.ENDS vias_gen$18$2$2$1$1$2

.SUBCKT nfet$2$2$2$1$1$2
.ENDS nfet$2$2$2$1$1$2

.SUBCKT vias_gen$7$2$2$1$1$2
.ENDS vias_gen$7$2$2$1$1$2

.SUBCKT vias_gen$10$1$1$2$1$1$2
.ENDS vias_gen$10$1$1$2$1$1$2

.SUBCKT vias_gen$2$1$1$1$2$1$1$2
.ENDS vias_gen$2$1$1$1$2$1$1$2

.SUBCKT pfet$2$1$1$2$1$1$2
.ENDS pfet$2$1$1$2$1$1$2

.SUBCKT vias_gen$6$1$1$2$1$1$2
.ENDS vias_gen$6$1$1$2$1$1$2

.SUBCKT vias_gen$18$1$1$2$1$1$2
.ENDS vias_gen$18$1$1$2$1$1$2

.SUBCKT nfet$2$1$1$2$1$1$2
.ENDS nfet$2$1$1$2$1$1$2

.SUBCKT vias_gen$7$1$1$2$1$1$2
.ENDS vias_gen$7$1$1$2$1$1$2

.SUBCKT vias_gen$10$2$1$2$1$2
.ENDS vias_gen$10$2$1$2$1$2

.SUBCKT vias_gen$2$1$2$1$2$1$2
.ENDS vias_gen$2$1$2$1$2$1$2

.SUBCKT pfet$2$2$1$2$1$2
.ENDS pfet$2$2$1$2$1$2

.SUBCKT vias_gen$6$2$1$2$1$2
.ENDS vias_gen$6$2$1$2$1$2

.SUBCKT vias_gen$18$2$1$2$1$2
.ENDS vias_gen$18$2$1$2$1$2

.SUBCKT nfet$2$2$1$2$1$2
.ENDS nfet$2$2$1$2$1$2

.SUBCKT vias_gen$7$2$1$2$1$2
.ENDS vias_gen$7$2$1$2$1$2

.SUBCKT vias_gen$10$1$1$1$2$1$2
.ENDS vias_gen$10$1$1$1$2$1$2

.SUBCKT vias_gen$2$1$1$1$1$2$1$2
.ENDS vias_gen$2$1$1$1$1$2$1$2

.SUBCKT pfet$2$1$1$1$2$1$2
.ENDS pfet$2$1$1$1$2$1$2

.SUBCKT vias_gen$6$1$1$1$2$1$2
.ENDS vias_gen$6$1$1$1$2$1$2

.SUBCKT vias_gen$18$1$1$1$2$1$2
.ENDS vias_gen$18$1$1$1$2$1$2

.SUBCKT nfet$2$1$1$1$2$1$2
.ENDS nfet$2$1$1$1$2$1$2

.SUBCKT vias_gen$7$1$1$1$2$1$2
.ENDS vias_gen$7$1$1$1$2$1$2

.SUBCKT vias_gen$10$3$2$1$2
.ENDS vias_gen$10$3$2$1$2

.SUBCKT vias_gen$2$1$3$2$1$2
.ENDS vias_gen$2$1$3$2$1$2

.SUBCKT pfet$2$3$2$1$2
.ENDS pfet$2$3$2$1$2

.SUBCKT vias_gen$6$3$2$1$2
.ENDS vias_gen$6$3$2$1$2

.SUBCKT vias_gen$18$3$2$1$2
.ENDS vias_gen$18$3$2$1$2

.SUBCKT nfet$2$3$2$1$2
.ENDS nfet$2$3$2$1$2

.SUBCKT vias_gen$7$3$2$1$2
.ENDS vias_gen$7$3$2$1$2

.SUBCKT vias_gen$10$1$2$2$1$2
.ENDS vias_gen$10$1$2$2$1$2

.SUBCKT vias_gen$2$1$1$2$2$1$2
.ENDS vias_gen$2$1$1$2$2$1$2

.SUBCKT pfet$2$1$2$2$1$2
.ENDS pfet$2$1$2$2$1$2

.SUBCKT vias_gen$6$1$2$2$1$2
.ENDS vias_gen$6$1$2$2$1$2

.SUBCKT vias_gen$18$1$2$2$1$2
.ENDS vias_gen$18$1$2$2$1$2

.SUBCKT nfet$2$1$2$2$1$2
.ENDS nfet$2$1$2$2$1$2

.SUBCKT vias_gen$7$1$2$2$1$2
.ENDS vias_gen$7$1$2$2$1$2

.SUBCKT vias_gen$10$2$1$1$1$3
.ENDS vias_gen$10$2$1$1$1$3

.SUBCKT vias_gen$2$1$2$1$1$1$3
.ENDS vias_gen$2$1$2$1$1$1$3

.SUBCKT pfet$2$2$1$1$1$3
.ENDS pfet$2$2$1$1$1$3

.SUBCKT vias_gen$6$2$1$1$1$3
.ENDS vias_gen$6$2$1$1$1$3

.SUBCKT vias_gen$18$2$1$1$1$3
.ENDS vias_gen$18$2$1$1$1$3

.SUBCKT nfet$2$2$1$1$1$3
.ENDS nfet$2$2$1$1$1$3

.SUBCKT vias_gen$7$2$1$1$1$3
.ENDS vias_gen$7$2$1$1$1$3

.SUBCKT vias_gen$10$1$1$1$1$1$3
.ENDS vias_gen$10$1$1$1$1$1$3

.SUBCKT vias_gen$2$1$1$1$1$1$1$3
.ENDS vias_gen$2$1$1$1$1$1$1$3

.SUBCKT pfet$2$1$1$1$1$1$3
.ENDS pfet$2$1$1$1$1$1$3

.SUBCKT vias_gen$6$1$1$1$1$1$3
.ENDS vias_gen$6$1$1$1$1$1$3

.SUBCKT vias_gen$18$1$1$1$1$1$3
.ENDS vias_gen$18$1$1$1$1$1$3

.SUBCKT nfet$2$1$1$1$1$1$3
.ENDS nfet$2$1$1$1$1$1$3

.SUBCKT vias_gen$7$1$1$1$1$1$3
.ENDS vias_gen$7$1$1$1$1$1$3

.SUBCKT vias_gen$10$3$1$1$3
.ENDS vias_gen$10$3$1$1$3

.SUBCKT vias_gen$2$1$3$1$1$3
.ENDS vias_gen$2$1$3$1$1$3

.SUBCKT pfet$2$3$1$1$3
.ENDS pfet$2$3$1$1$3

.SUBCKT vias_gen$6$3$1$1$3
.ENDS vias_gen$6$3$1$1$3

.SUBCKT vias_gen$18$3$1$1$3
.ENDS vias_gen$18$3$1$1$3

.SUBCKT nfet$2$3$1$1$3
.ENDS nfet$2$3$1$1$3

.SUBCKT vias_gen$7$3$1$1$3
.ENDS vias_gen$7$3$1$1$3

.SUBCKT vias_gen$10$1$2$1$1$3
.ENDS vias_gen$10$1$2$1$1$3

.SUBCKT vias_gen$2$1$1$2$1$1$3
.ENDS vias_gen$2$1$1$2$1$1$3

.SUBCKT pfet$2$1$2$1$1$3
.ENDS pfet$2$1$2$1$1$3

.SUBCKT vias_gen$6$1$2$1$1$3
.ENDS vias_gen$6$1$2$1$1$3

.SUBCKT vias_gen$18$1$2$1$1$3
.ENDS vias_gen$18$1$2$1$1$3

.SUBCKT nfet$2$1$2$1$1$3
.ENDS nfet$2$1$2$1$1$3

.SUBCKT vias_gen$7$1$2$1$1$3
.ENDS vias_gen$7$1$2$1$1$3

.SUBCKT vias_gen$10$2$1$1$1$1$1
.ENDS vias_gen$10$2$1$1$1$1$1

.SUBCKT vias_gen$2$1$2$1$1$1$1$1
.ENDS vias_gen$2$1$2$1$1$1$1$1

.SUBCKT pfet$2$2$1$1$1$1$1
.ENDS pfet$2$2$1$1$1$1$1

.SUBCKT vias_gen$6$2$1$1$1$1$1
.ENDS vias_gen$6$2$1$1$1$1$1

.SUBCKT vias_gen$18$2$1$1$1$1$1
.ENDS vias_gen$18$2$1$1$1$1$1

.SUBCKT nfet$2$2$1$1$1$1$1
.ENDS nfet$2$2$1$1$1$1$1

.SUBCKT vias_gen$7$2$1$1$1$1$1
.ENDS vias_gen$7$2$1$1$1$1$1

.SUBCKT vias_gen$10$1$1$1$1$1$1$1
.ENDS vias_gen$10$1$1$1$1$1$1$1

.SUBCKT vias_gen$2$1$1$1$1$1$1$1$1
.ENDS vias_gen$2$1$1$1$1$1$1$1$1

.SUBCKT pfet$2$1$1$1$1$1$1$1
.ENDS pfet$2$1$1$1$1$1$1$1

.SUBCKT vias_gen$6$1$1$1$1$1$1$1
.ENDS vias_gen$6$1$1$1$1$1$1$1

.SUBCKT vias_gen$18$1$1$1$1$1$1$1
.ENDS vias_gen$18$1$1$1$1$1$1$1

.SUBCKT nfet$2$1$1$1$1$1$1$1
.ENDS nfet$2$1$1$1$1$1$1$1

.SUBCKT vias_gen$7$1$1$1$1$1$1$1
.ENDS vias_gen$7$1$1$1$1$1$1$1

.SUBCKT vias_gen$10$3$1$1$1$1
.ENDS vias_gen$10$3$1$1$1$1

.SUBCKT vias_gen$2$1$3$1$1$1$1
.ENDS vias_gen$2$1$3$1$1$1$1

.SUBCKT pfet$2$3$1$1$1$1
.ENDS pfet$2$3$1$1$1$1

.SUBCKT vias_gen$6$3$1$1$1$1
.ENDS vias_gen$6$3$1$1$1$1

.SUBCKT vias_gen$18$3$1$1$1$1
.ENDS vias_gen$18$3$1$1$1$1

.SUBCKT nfet$2$3$1$1$1$1
.ENDS nfet$2$3$1$1$1$1

.SUBCKT vias_gen$7$3$1$1$1$1
.ENDS vias_gen$7$3$1$1$1$1

.SUBCKT vias_gen$10$1$2$1$1$1$1
.ENDS vias_gen$10$1$2$1$1$1$1

.SUBCKT vias_gen$2$1$1$2$1$1$1$1
.ENDS vias_gen$2$1$1$2$1$1$1$1

.SUBCKT pfet$2$1$2$1$1$1$1
.ENDS pfet$2$1$2$1$1$1$1

.SUBCKT vias_gen$6$1$2$1$1$1$1
.ENDS vias_gen$6$1$2$1$1$1$1

.SUBCKT vias_gen$18$1$2$1$1$1$1
.ENDS vias_gen$18$1$2$1$1$1$1

.SUBCKT nfet$2$1$2$1$1$1$1
.ENDS nfet$2$1$2$1$1$1$1

.SUBCKT vias_gen$7$1$2$1$1$1$1
.ENDS vias_gen$7$1$2$1$1$1$1

.SUBCKT vias_gen$10$2$2$1$1$1
.ENDS vias_gen$10$2$2$1$1$1

.SUBCKT vias_gen$2$1$2$2$1$1$1
.ENDS vias_gen$2$1$2$2$1$1$1

.SUBCKT pfet$2$2$2$1$1$1
.ENDS pfet$2$2$2$1$1$1

.SUBCKT vias_gen$6$2$2$1$1$1
.ENDS vias_gen$6$2$2$1$1$1

.SUBCKT vias_gen$18$2$2$1$1$1
.ENDS vias_gen$18$2$2$1$1$1

.SUBCKT nfet$2$2$2$1$1$1
.ENDS nfet$2$2$2$1$1$1

.SUBCKT vias_gen$7$2$2$1$1$1
.ENDS vias_gen$7$2$2$1$1$1

.SUBCKT vias_gen$10$1$1$2$1$1$1
.ENDS vias_gen$10$1$1$2$1$1$1

.SUBCKT vias_gen$2$1$1$1$2$1$1$1
.ENDS vias_gen$2$1$1$1$2$1$1$1

.SUBCKT pfet$2$1$1$2$1$1$1
.ENDS pfet$2$1$1$2$1$1$1

.SUBCKT vias_gen$6$1$1$2$1$1$1
.ENDS vias_gen$6$1$1$2$1$1$1

.SUBCKT vias_gen$18$1$1$2$1$1$1
.ENDS vias_gen$18$1$1$2$1$1$1

.SUBCKT nfet$2$1$1$2$1$1$1
.ENDS nfet$2$1$1$2$1$1$1

.SUBCKT vias_gen$7$1$1$2$1$1$1
.ENDS vias_gen$7$1$1$2$1$1$1

.SUBCKT vias_gen$10$2$1$2$1$1
.ENDS vias_gen$10$2$1$2$1$1

.SUBCKT vias_gen$2$1$2$1$2$1$1
.ENDS vias_gen$2$1$2$1$2$1$1

.SUBCKT pfet$2$2$1$2$1$1
.ENDS pfet$2$2$1$2$1$1

.SUBCKT vias_gen$6$2$1$2$1$1
.ENDS vias_gen$6$2$1$2$1$1

.SUBCKT vias_gen$18$2$1$2$1$1
.ENDS vias_gen$18$2$1$2$1$1

.SUBCKT nfet$2$2$1$2$1$1
.ENDS nfet$2$2$1$2$1$1

.SUBCKT vias_gen$7$2$1$2$1$1
.ENDS vias_gen$7$2$1$2$1$1

.SUBCKT vias_gen$10$1$1$1$2$1$1
.ENDS vias_gen$10$1$1$1$2$1$1

.SUBCKT vias_gen$2$1$1$1$1$2$1$1
.ENDS vias_gen$2$1$1$1$1$2$1$1

.SUBCKT pfet$2$1$1$1$2$1$1
.ENDS pfet$2$1$1$1$2$1$1

.SUBCKT vias_gen$6$1$1$1$2$1$1
.ENDS vias_gen$6$1$1$1$2$1$1

.SUBCKT vias_gen$18$1$1$1$2$1$1
.ENDS vias_gen$18$1$1$1$2$1$1

.SUBCKT nfet$2$1$1$1$2$1$1
.ENDS nfet$2$1$1$1$2$1$1

.SUBCKT vias_gen$7$1$1$1$2$1$1
.ENDS vias_gen$7$1$1$1$2$1$1

.SUBCKT vias_gen$10$3$2$1$1
.ENDS vias_gen$10$3$2$1$1

.SUBCKT vias_gen$2$1$3$2$1$1
.ENDS vias_gen$2$1$3$2$1$1

.SUBCKT pfet$2$3$2$1$1
.ENDS pfet$2$3$2$1$1

.SUBCKT vias_gen$6$3$2$1$1
.ENDS vias_gen$6$3$2$1$1

.SUBCKT vias_gen$18$3$2$1$1
.ENDS vias_gen$18$3$2$1$1

.SUBCKT nfet$2$3$2$1$1
.ENDS nfet$2$3$2$1$1

.SUBCKT vias_gen$7$3$2$1$1
.ENDS vias_gen$7$3$2$1$1

.SUBCKT vias_gen$10$1$2$2$1$1
.ENDS vias_gen$10$1$2$2$1$1

.SUBCKT vias_gen$2$1$1$2$2$1$1
.ENDS vias_gen$2$1$1$2$2$1$1

.SUBCKT pfet$2$1$2$2$1$1
.ENDS pfet$2$1$2$2$1$1

.SUBCKT vias_gen$6$1$2$2$1$1
.ENDS vias_gen$6$1$2$2$1$1

.SUBCKT vias_gen$18$1$2$2$1$1
.ENDS vias_gen$18$1$2$2$1$1

.SUBCKT nfet$2$1$2$2$1$1
.ENDS nfet$2$1$2$2$1$1

.SUBCKT vias_gen$7$1$2$2$1$1
.ENDS vias_gen$7$1$2$2$1$1

.SUBCKT vias_gen$10$2$1$1$1$2
.ENDS vias_gen$10$2$1$1$1$2

.SUBCKT vias_gen$2$1$2$1$1$1$2
.ENDS vias_gen$2$1$2$1$1$1$2

.SUBCKT pfet$2$2$1$1$1$2
.ENDS pfet$2$2$1$1$1$2

.SUBCKT vias_gen$6$2$1$1$1$2
.ENDS vias_gen$6$2$1$1$1$2

.SUBCKT vias_gen$18$2$1$1$1$2
.ENDS vias_gen$18$2$1$1$1$2

.SUBCKT nfet$2$2$1$1$1$2
.ENDS nfet$2$2$1$1$1$2

.SUBCKT vias_gen$7$2$1$1$1$2
.ENDS vias_gen$7$2$1$1$1$2

.SUBCKT vias_gen$10$1$1$1$1$1$2
.ENDS vias_gen$10$1$1$1$1$1$2

.SUBCKT vias_gen$2$1$1$1$1$1$1$2
.ENDS vias_gen$2$1$1$1$1$1$1$2

.SUBCKT pfet$2$1$1$1$1$1$2
.ENDS pfet$2$1$1$1$1$1$2

.SUBCKT vias_gen$6$1$1$1$1$1$2
.ENDS vias_gen$6$1$1$1$1$1$2

.SUBCKT vias_gen$18$1$1$1$1$1$2
.ENDS vias_gen$18$1$1$1$1$1$2

.SUBCKT nfet$2$1$1$1$1$1$2
.ENDS nfet$2$1$1$1$1$1$2

.SUBCKT vias_gen$7$1$1$1$1$1$2
.ENDS vias_gen$7$1$1$1$1$1$2

.SUBCKT vias_gen$10$3$1$1$2
.ENDS vias_gen$10$3$1$1$2

.SUBCKT vias_gen$2$1$3$1$1$2
.ENDS vias_gen$2$1$3$1$1$2

.SUBCKT pfet$2$3$1$1$2
.ENDS pfet$2$3$1$1$2

.SUBCKT vias_gen$6$3$1$1$2
.ENDS vias_gen$6$3$1$1$2

.SUBCKT vias_gen$18$3$1$1$2
.ENDS vias_gen$18$3$1$1$2

.SUBCKT nfet$2$3$1$1$2
.ENDS nfet$2$3$1$1$2

.SUBCKT vias_gen$7$3$1$1$2
.ENDS vias_gen$7$3$1$1$2

.SUBCKT vias_gen$10$1$2$1$1$2
.ENDS vias_gen$10$1$2$1$1$2

.SUBCKT vias_gen$2$1$1$2$1$1$2
.ENDS vias_gen$2$1$1$2$1$1$2

.SUBCKT pfet$2$1$2$1$1$2
.ENDS pfet$2$1$2$1$1$2

.SUBCKT vias_gen$6$1$2$1$1$2
.ENDS vias_gen$6$1$2$1$1$2

.SUBCKT vias_gen$18$1$2$1$1$2
.ENDS vias_gen$18$1$2$1$1$2

.SUBCKT nfet$2$1$2$1$1$2
.ENDS nfet$2$1$2$1$1$2

.SUBCKT vias_gen$7$1$2$1$1$2
.ENDS vias_gen$7$1$2$1$1$2

.SUBCKT vias_gen$10$2$2$1$2
.ENDS vias_gen$10$2$2$1$2

.SUBCKT vias_gen$2$1$2$2$1$2
.ENDS vias_gen$2$1$2$2$1$2

.SUBCKT pfet$2$2$2$1$2
.ENDS pfet$2$2$2$1$2

.SUBCKT vias_gen$6$2$2$1$2
.ENDS vias_gen$6$2$2$1$2

.SUBCKT vias_gen$18$2$2$1$2
.ENDS vias_gen$18$2$2$1$2

.SUBCKT nfet$2$2$2$1$2
.ENDS nfet$2$2$2$1$2

.SUBCKT vias_gen$7$2$2$1$2
.ENDS vias_gen$7$2$2$1$2

.SUBCKT vias_gen$10$1$1$2$1$2
.ENDS vias_gen$10$1$1$2$1$2

.SUBCKT vias_gen$2$1$1$1$2$1$2
.ENDS vias_gen$2$1$1$1$2$1$2

.SUBCKT pfet$2$1$1$2$1$2
.ENDS pfet$2$1$1$2$1$2

.SUBCKT vias_gen$6$1$1$2$1$2
.ENDS vias_gen$6$1$1$2$1$2

.SUBCKT vias_gen$18$1$1$2$1$2
.ENDS vias_gen$18$1$1$2$1$2

.SUBCKT nfet$2$1$1$2$1$2
.ENDS nfet$2$1$1$2$1$2

.SUBCKT vias_gen$7$1$1$2$1$2
.ENDS vias_gen$7$1$1$2$1$2

.SUBCKT vias_gen$10$2$1$2$2
.ENDS vias_gen$10$2$1$2$2

.SUBCKT vias_gen$2$1$2$1$2$2
.ENDS vias_gen$2$1$2$1$2$2

.SUBCKT pfet$2$2$1$2$2
.ENDS pfet$2$2$1$2$2

.SUBCKT vias_gen$6$2$1$2$2
.ENDS vias_gen$6$2$1$2$2

.SUBCKT vias_gen$18$2$1$2$2
.ENDS vias_gen$18$2$1$2$2

.SUBCKT nfet$2$2$1$2$2
.ENDS nfet$2$2$1$2$2

.SUBCKT vias_gen$7$2$1$2$2
.ENDS vias_gen$7$2$1$2$2

.SUBCKT vias_gen$10$1$1$1$2$2
.ENDS vias_gen$10$1$1$1$2$2

.SUBCKT vias_gen$2$1$1$1$1$2$2
.ENDS vias_gen$2$1$1$1$1$2$2

.SUBCKT pfet$2$1$1$1$2$2
.ENDS pfet$2$1$1$1$2$2

.SUBCKT vias_gen$6$1$1$1$2$2
.ENDS vias_gen$6$1$1$1$2$2

.SUBCKT vias_gen$18$1$1$1$2$2
.ENDS vias_gen$18$1$1$1$2$2

.SUBCKT nfet$2$1$1$1$2$2
.ENDS nfet$2$1$1$1$2$2

.SUBCKT vias_gen$7$1$1$1$2$2
.ENDS vias_gen$7$1$1$1$2$2

.SUBCKT vias_gen$10$3$2$2
.ENDS vias_gen$10$3$2$2

.SUBCKT vias_gen$2$1$3$2$2
.ENDS vias_gen$2$1$3$2$2

.SUBCKT pfet$2$3$2$2
.ENDS pfet$2$3$2$2

.SUBCKT vias_gen$6$3$2$2
.ENDS vias_gen$6$3$2$2

.SUBCKT vias_gen$18$3$2$2
.ENDS vias_gen$18$3$2$2

.SUBCKT nfet$2$3$2$2
.ENDS nfet$2$3$2$2

.SUBCKT vias_gen$7$3$2$2
.ENDS vias_gen$7$3$2$2

.SUBCKT vias_gen$10$1$2$2$2
.ENDS vias_gen$10$1$2$2$2

.SUBCKT vias_gen$2$1$1$2$2$2
.ENDS vias_gen$2$1$1$2$2$2

.SUBCKT pfet$2$1$2$2$2
.ENDS pfet$2$1$2$2$2

.SUBCKT vias_gen$6$1$2$2$2
.ENDS vias_gen$6$1$2$2$2

.SUBCKT vias_gen$18$1$2$2$2
.ENDS vias_gen$18$1$2$2$2

.SUBCKT nfet$2$1$2$2$2
.ENDS nfet$2$1$2$2$2

.SUBCKT vias_gen$7$1$2$2$2
.ENDS vias_gen$7$1$2$2$2

.SUBCKT vias_gen$10$3$1$1$1
.ENDS vias_gen$10$3$1$1$1

.SUBCKT vias_gen$2$1$3$1$1$1
.ENDS vias_gen$2$1$3$1$1$1

.SUBCKT pfet$2$3$1$1$1
.ENDS pfet$2$3$1$1$1

.SUBCKT vias_gen$6$3$1$1$1
.ENDS vias_gen$6$3$1$1$1

.SUBCKT vias_gen$18$3$1$1$1
.ENDS vias_gen$18$3$1$1$1

.SUBCKT nfet$2$3$1$1$1
.ENDS nfet$2$3$1$1$1

.SUBCKT vias_gen$7$3$1$1$1
.ENDS vias_gen$7$3$1$1$1

.SUBCKT vias_gen$10$1$2$1$1$1
.ENDS vias_gen$10$1$2$1$1$1

.SUBCKT vias_gen$2$1$1$2$1$1$1
.ENDS vias_gen$2$1$1$2$1$1$1

.SUBCKT pfet$2$1$2$1$1$1
.ENDS pfet$2$1$2$1$1$1

.SUBCKT vias_gen$6$1$2$1$1$1
.ENDS vias_gen$6$1$2$1$1$1

.SUBCKT vias_gen$18$1$2$1$1$1
.ENDS vias_gen$18$1$2$1$1$1

.SUBCKT nfet$2$1$2$1$1$1
.ENDS nfet$2$1$2$1$1$1

.SUBCKT vias_gen$7$1$2$1$1$1
.ENDS vias_gen$7$1$2$1$1$1

.SUBCKT vias_gen$10$2$2$1$1
.ENDS vias_gen$10$2$2$1$1

.SUBCKT vias_gen$2$1$2$2$1$1
.ENDS vias_gen$2$1$2$2$1$1

.SUBCKT pfet$2$2$2$1$1
.ENDS pfet$2$2$2$1$1

.SUBCKT vias_gen$6$2$2$1$1
.ENDS vias_gen$6$2$2$1$1

.SUBCKT vias_gen$18$2$2$1$1
.ENDS vias_gen$18$2$2$1$1

.SUBCKT nfet$2$2$2$1$1
.ENDS nfet$2$2$2$1$1

.SUBCKT vias_gen$7$2$2$1$1
.ENDS vias_gen$7$2$2$1$1

.SUBCKT vias_gen$10$1$1$2$1$1
.ENDS vias_gen$10$1$1$2$1$1

.SUBCKT vias_gen$2$1$1$1$2$1$1
.ENDS vias_gen$2$1$1$1$2$1$1

.SUBCKT pfet$2$1$1$2$1$1
.ENDS pfet$2$1$1$2$1$1

.SUBCKT vias_gen$6$1$1$2$1$1
.ENDS vias_gen$6$1$1$2$1$1

.SUBCKT vias_gen$18$1$1$2$1$1
.ENDS vias_gen$18$1$1$2$1$1

.SUBCKT nfet$2$1$1$2$1$1
.ENDS nfet$2$1$1$2$1$1

.SUBCKT vias_gen$7$1$1$2$1$1
.ENDS vias_gen$7$1$1$2$1$1

.SUBCKT vias_gen$10$2$1$2$1
.ENDS vias_gen$10$2$1$2$1

.SUBCKT vias_gen$2$1$2$1$2$1
.ENDS vias_gen$2$1$2$1$2$1

.SUBCKT pfet$2$2$1$2$1
.ENDS pfet$2$2$1$2$1

.SUBCKT vias_gen$6$2$1$2$1
.ENDS vias_gen$6$2$1$2$1

.SUBCKT vias_gen$18$2$1$2$1
.ENDS vias_gen$18$2$1$2$1

.SUBCKT nfet$2$2$1$2$1
.ENDS nfet$2$2$1$2$1

.SUBCKT vias_gen$7$2$1$2$1
.ENDS vias_gen$7$2$1$2$1

.SUBCKT vias_gen$10$1$1$1$2$1
.ENDS vias_gen$10$1$1$1$2$1

.SUBCKT vias_gen$2$1$1$1$1$2$1
.ENDS vias_gen$2$1$1$1$1$2$1

.SUBCKT pfet$2$1$1$1$2$1
.ENDS pfet$2$1$1$1$2$1

.SUBCKT vias_gen$6$1$1$1$2$1
.ENDS vias_gen$6$1$1$1$2$1

.SUBCKT vias_gen$18$1$1$1$2$1
.ENDS vias_gen$18$1$1$1$2$1

.SUBCKT nfet$2$1$1$1$2$1
.ENDS nfet$2$1$1$1$2$1

.SUBCKT vias_gen$7$1$1$1$2$1
.ENDS vias_gen$7$1$1$1$2$1

.SUBCKT vias_gen$10$3$2$1
.ENDS vias_gen$10$3$2$1

.SUBCKT vias_gen$2$1$3$2$1
.ENDS vias_gen$2$1$3$2$1

.SUBCKT pfet$2$3$2$1
.ENDS pfet$2$3$2$1

.SUBCKT vias_gen$6$3$2$1
.ENDS vias_gen$6$3$2$1

.SUBCKT vias_gen$18$3$2$1
.ENDS vias_gen$18$3$2$1

.SUBCKT nfet$2$3$2$1
.ENDS nfet$2$3$2$1

.SUBCKT vias_gen$7$3$2$1
.ENDS vias_gen$7$3$2$1

.SUBCKT vias_gen$10$1$2$2$1
.ENDS vias_gen$10$1$2$2$1

.SUBCKT vias_gen$2$1$1$2$2$1
.ENDS vias_gen$2$1$1$2$2$1

.SUBCKT pfet$2$1$2$2$1
.ENDS pfet$2$1$2$2$1

.SUBCKT vias_gen$6$1$2$2$1
.ENDS vias_gen$6$1$2$2$1

.SUBCKT vias_gen$18$1$2$2$1
.ENDS vias_gen$18$1$2$2$1

.SUBCKT nfet$2$1$2$2$1
.ENDS nfet$2$1$2$2$1

.SUBCKT vias_gen$7$1$2$2$1
.ENDS vias_gen$7$1$2$2$1

.SUBCKT vias_gen$10$2$1$1$1
.ENDS vias_gen$10$2$1$1$1

.SUBCKT vias_gen$2$1$2$1$1$1
.ENDS vias_gen$2$1$2$1$1$1

.SUBCKT pfet$2$2$1$1$1
.ENDS pfet$2$2$1$1$1

.SUBCKT vias_gen$6$2$1$1$1
.ENDS vias_gen$6$2$1$1$1

.SUBCKT vias_gen$18$2$1$1$1
.ENDS vias_gen$18$2$1$1$1

.SUBCKT nfet$2$2$1$1$1
.ENDS nfet$2$2$1$1$1

.SUBCKT vias_gen$7$2$1$1$1
.ENDS vias_gen$7$2$1$1$1

.SUBCKT vias_gen$10$1$1$1$1$1
.ENDS vias_gen$10$1$1$1$1$1

.SUBCKT vias_gen$2$1$1$1$1$1$1
.ENDS vias_gen$2$1$1$1$1$1$1

.SUBCKT pfet$2$1$1$1$1$1
.ENDS pfet$2$1$1$1$1$1

.SUBCKT vias_gen$6$1$1$1$1$1
.ENDS vias_gen$6$1$1$1$1$1

.SUBCKT vias_gen$18$1$1$1$1$1
.ENDS vias_gen$18$1$1$1$1$1

.SUBCKT nfet$2$1$1$1$1$1
.ENDS nfet$2$1$1$1$1$1

.SUBCKT vias_gen$7$1$1$1$1$1
.ENDS vias_gen$7$1$1$1$1$1

.SUBCKT vias_gen$10$3$1$1
.ENDS vias_gen$10$3$1$1

.SUBCKT vias_gen$2$1$3$1$1
.ENDS vias_gen$2$1$3$1$1

.SUBCKT pfet$2$3$1$1
.ENDS pfet$2$3$1$1

.SUBCKT vias_gen$6$3$1$1
.ENDS vias_gen$6$3$1$1

.SUBCKT vias_gen$18$3$1$1
.ENDS vias_gen$18$3$1$1

.SUBCKT nfet$2$3$1$1
.ENDS nfet$2$3$1$1

.SUBCKT vias_gen$7$3$1$1
.ENDS vias_gen$7$3$1$1

.SUBCKT vias_gen$10$1$2$1$1
.ENDS vias_gen$10$1$2$1$1

.SUBCKT vias_gen$2$1$1$2$1$1
.ENDS vias_gen$2$1$1$2$1$1

.SUBCKT pfet$2$1$2$1$1
.ENDS pfet$2$1$2$1$1

.SUBCKT vias_gen$6$1$2$1$1
.ENDS vias_gen$6$1$2$1$1

.SUBCKT vias_gen$18$1$2$1$1
.ENDS vias_gen$18$1$2$1$1

.SUBCKT nfet$2$1$2$1$1
.ENDS nfet$2$1$2$1$1

.SUBCKT vias_gen$7$1$2$1$1
.ENDS vias_gen$7$1$2$1$1

.SUBCKT vias_gen$10$2$2$1
.ENDS vias_gen$10$2$2$1

.SUBCKT vias_gen$2$1$2$2$1
.ENDS vias_gen$2$1$2$2$1

.SUBCKT pfet$2$2$2$1
.ENDS pfet$2$2$2$1

.SUBCKT vias_gen$6$2$2$1
.ENDS vias_gen$6$2$2$1

.SUBCKT vias_gen$18$2$2$1
.ENDS vias_gen$18$2$2$1

.SUBCKT nfet$2$2$2$1
.ENDS nfet$2$2$2$1

.SUBCKT vias_gen$7$2$2$1
.ENDS vias_gen$7$2$2$1

.SUBCKT vias_gen$10$1$1$2$1
.ENDS vias_gen$10$1$1$2$1

.SUBCKT vias_gen$2$1$1$1$2$1
.ENDS vias_gen$2$1$1$1$2$1

.SUBCKT pfet$2$1$1$2$1
.ENDS pfet$2$1$1$2$1

.SUBCKT vias_gen$6$1$1$2$1
.ENDS vias_gen$6$1$1$2$1

.SUBCKT vias_gen$18$1$1$2$1
.ENDS vias_gen$18$1$1$2$1

.SUBCKT nfet$2$1$1$2$1
.ENDS nfet$2$1$1$2$1

.SUBCKT vias_gen$7$1$1$2$1
.ENDS vias_gen$7$1$1$2$1

.SUBCKT vias_gen$10$2$1$2
.ENDS vias_gen$10$2$1$2

.SUBCKT vias_gen$2$1$2$1$2
.ENDS vias_gen$2$1$2$1$2

.SUBCKT pfet$2$2$1$2
.ENDS pfet$2$2$1$2

.SUBCKT vias_gen$6$2$1$2
.ENDS vias_gen$6$2$1$2

.SUBCKT vias_gen$18$2$1$2
.ENDS vias_gen$18$2$1$2

.SUBCKT nfet$2$2$1$2
.ENDS nfet$2$2$1$2

.SUBCKT vias_gen$7$2$1$2
.ENDS vias_gen$7$2$1$2

.SUBCKT vias_gen$10$1$1$1$2
.ENDS vias_gen$10$1$1$1$2

.SUBCKT vias_gen$2$1$1$1$1$2
.ENDS vias_gen$2$1$1$1$1$2

.SUBCKT pfet$2$1$1$1$2
.ENDS pfet$2$1$1$1$2

.SUBCKT vias_gen$6$1$1$1$2
.ENDS vias_gen$6$1$1$1$2

.SUBCKT vias_gen$18$1$1$1$2
.ENDS vias_gen$18$1$1$1$2

.SUBCKT nfet$2$1$1$1$2
.ENDS nfet$2$1$1$1$2

.SUBCKT vias_gen$7$1$1$1$2
.ENDS vias_gen$7$1$1$1$2

.SUBCKT vias_gen$10$3$2
.ENDS vias_gen$10$3$2

.SUBCKT vias_gen$2$1$3$2
.ENDS vias_gen$2$1$3$2

.SUBCKT pfet$2$3$2
.ENDS pfet$2$3$2

.SUBCKT vias_gen$6$3$2
.ENDS vias_gen$6$3$2

.SUBCKT vias_gen$18$3$2
.ENDS vias_gen$18$3$2

.SUBCKT nfet$2$3$2
.ENDS nfet$2$3$2

.SUBCKT vias_gen$7$3$2
.ENDS vias_gen$7$3$2

.SUBCKT vias_gen$10$1$2$2
.ENDS vias_gen$10$1$2$2

.SUBCKT vias_gen$2$1$1$2$2
.ENDS vias_gen$2$1$1$2$2

.SUBCKT pfet$2$1$2$2
.ENDS pfet$2$1$2$2

.SUBCKT vias_gen$6$1$2$2
.ENDS vias_gen$6$1$2$2

.SUBCKT vias_gen$18$1$2$2
.ENDS vias_gen$18$1$2$2

.SUBCKT nfet$2$1$2$2
.ENDS nfet$2$1$2$2

.SUBCKT vias_gen$7$1$2$2
.ENDS vias_gen$7$1$2$2

.SUBCKT vias_gen$10$2$1$1
.ENDS vias_gen$10$2$1$1

.SUBCKT vias_gen$2$1$2$1$1
.ENDS vias_gen$2$1$2$1$1

.SUBCKT pfet$2$2$1$1
.ENDS pfet$2$2$1$1

.SUBCKT vias_gen$6$2$1$1
.ENDS vias_gen$6$2$1$1

.SUBCKT vias_gen$18$2$1$1
.ENDS vias_gen$18$2$1$1

.SUBCKT nfet$2$2$1$1
.ENDS nfet$2$2$1$1

.SUBCKT vias_gen$7$2$1$1
.ENDS vias_gen$7$2$1$1

.SUBCKT vias_gen$10$1$1$1$1
.ENDS vias_gen$10$1$1$1$1

.SUBCKT vias_gen$2$1$1$1$1$1
.ENDS vias_gen$2$1$1$1$1$1

.SUBCKT pfet$2$1$1$1$1
.ENDS pfet$2$1$1$1$1

.SUBCKT vias_gen$6$1$1$1$1
.ENDS vias_gen$6$1$1$1$1

.SUBCKT vias_gen$18$1$1$1$1
.ENDS vias_gen$18$1$1$1$1

.SUBCKT nfet$2$1$1$1$1
.ENDS nfet$2$1$1$1$1

.SUBCKT vias_gen$7$1$1$1$1
.ENDS vias_gen$7$1$1$1$1

.SUBCKT vias_gen$10$3$1
.ENDS vias_gen$10$3$1

.SUBCKT vias_gen$2$1$3$1
.ENDS vias_gen$2$1$3$1

.SUBCKT pfet$2$3$1
.ENDS pfet$2$3$1

.SUBCKT vias_gen$6$3$1
.ENDS vias_gen$6$3$1

.SUBCKT vias_gen$18$3$1
.ENDS vias_gen$18$3$1

.SUBCKT nfet$2$3$1
.ENDS nfet$2$3$1

.SUBCKT vias_gen$7$3$1
.ENDS vias_gen$7$3$1

.SUBCKT vias_gen$10$1$2$1
.ENDS vias_gen$10$1$2$1

.SUBCKT vias_gen$2$1$1$2$1
.ENDS vias_gen$2$1$1$2$1

.SUBCKT pfet$2$1$2$1
.ENDS pfet$2$1$2$1

.SUBCKT vias_gen$6$1$2$1
.ENDS vias_gen$6$1$2$1

.SUBCKT vias_gen$18$1$2$1
.ENDS vias_gen$18$1$2$1

.SUBCKT nfet$2$1$2$1
.ENDS nfet$2$1$2$1

.SUBCKT vias_gen$7$1$2$1
.ENDS vias_gen$7$1$2$1

.SUBCKT vias_gen$10$2$2
.ENDS vias_gen$10$2$2

.SUBCKT vias_gen$2$1$2$2
.ENDS vias_gen$2$1$2$2

.SUBCKT pfet$2$2$2
.ENDS pfet$2$2$2

.SUBCKT vias_gen$6$2$2
.ENDS vias_gen$6$2$2

.SUBCKT vias_gen$18$2$2
.ENDS vias_gen$18$2$2

.SUBCKT nfet$2$2$2
.ENDS nfet$2$2$2

.SUBCKT vias_gen$7$2$2
.ENDS vias_gen$7$2$2

.SUBCKT vias_gen$10$1$1$2
.ENDS vias_gen$10$1$1$2

.SUBCKT vias_gen$2$1$1$1$2
.ENDS vias_gen$2$1$1$1$2

.SUBCKT pfet$2$1$1$2
.ENDS pfet$2$1$1$2

.SUBCKT vias_gen$6$1$1$2
.ENDS vias_gen$6$1$1$2

.SUBCKT vias_gen$18$1$1$2
.ENDS vias_gen$18$1$1$2

.SUBCKT nfet$2$1$1$2
.ENDS nfet$2$1$1$2

.SUBCKT vias_gen$7$1$1$2
.ENDS vias_gen$7$1$1$2

.SUBCKT vias_gen$10$2$1
.ENDS vias_gen$10$2$1

.SUBCKT vias_gen$2$1$2$1
.ENDS vias_gen$2$1$2$1

.SUBCKT pfet$2$2$1
.ENDS pfet$2$2$1

.SUBCKT vias_gen$6$2$1
.ENDS vias_gen$6$2$1

.SUBCKT vias_gen$18$2$1
.ENDS vias_gen$18$2$1

.SUBCKT nfet$2$2$1
.ENDS nfet$2$2$1

.SUBCKT vias_gen$7$2$1
.ENDS vias_gen$7$2$1

.SUBCKT vias_gen$10$1$1$1
.ENDS vias_gen$10$1$1$1

.SUBCKT vias_gen$2$1$1$1$1
.ENDS vias_gen$2$1$1$1$1

.SUBCKT pfet$2$1$1$1
.ENDS pfet$2$1$1$1

.SUBCKT vias_gen$6$1$1$1
.ENDS vias_gen$6$1$1$1

.SUBCKT vias_gen$18$1$1$1
.ENDS vias_gen$18$1$1$1

.SUBCKT nfet$2$1$1$1
.ENDS nfet$2$1$1$1

.SUBCKT vias_gen$7$1$1$1
.ENDS vias_gen$7$1$1$1

.SUBCKT vias_gen$10$3
.ENDS vias_gen$10$3

.SUBCKT vias_gen$2$1$3
.ENDS vias_gen$2$1$3

.SUBCKT pfet$2$3
.ENDS pfet$2$3

.SUBCKT vias_gen$6$3
.ENDS vias_gen$6$3

.SUBCKT vias_gen$18$3
.ENDS vias_gen$18$3

.SUBCKT nfet$2$3
.ENDS nfet$2$3

.SUBCKT vias_gen$7$3
.ENDS vias_gen$7$3

.SUBCKT vias_gen$10$1$2
.ENDS vias_gen$10$1$2

.SUBCKT vias_gen$2$1$1$2
.ENDS vias_gen$2$1$1$2

.SUBCKT pfet$2$1$2
.ENDS pfet$2$1$2

.SUBCKT vias_gen$6$1$2
.ENDS vias_gen$6$1$2

.SUBCKT vias_gen$18$1$2
.ENDS vias_gen$18$1$2

.SUBCKT nfet$2$1$2
.ENDS nfet$2$1$2

.SUBCKT vias_gen$7$1$2
.ENDS vias_gen$7$1$2

.SUBCKT vias_gen$10$2
.ENDS vias_gen$10$2

.SUBCKT vias_gen$2$1$2
.ENDS vias_gen$2$1$2

.SUBCKT pfet$2$2
.ENDS pfet$2$2

.SUBCKT vias_gen$6$2
.ENDS vias_gen$6$2

.SUBCKT vias_gen$18$2
.ENDS vias_gen$18$2

.SUBCKT nfet$2$2
.ENDS nfet$2$2

.SUBCKT vias_gen$7$2
.ENDS vias_gen$7$2

.SUBCKT vias_gen$10$1$1
.ENDS vias_gen$10$1$1

.SUBCKT vias_gen$2$1$1$1
.ENDS vias_gen$2$1$1$1

.SUBCKT pfet$2$1$1
.ENDS pfet$2$1$1

.SUBCKT vias_gen$6$1$1
.ENDS vias_gen$6$1$1

.SUBCKT vias_gen$18$1$1
.ENDS vias_gen$18$1$1

.SUBCKT nfet$2$1$1
.ENDS nfet$2$1$1

.SUBCKT vias_gen$7$1$1
.ENDS vias_gen$7$1$1

.SUBCKT vias_gen$10
.ENDS vias_gen$10

.SUBCKT vias_gen$2$1
.ENDS vias_gen$2$1

.SUBCKT pfet$2
.ENDS pfet$2

.SUBCKT vias_gen$6
.ENDS vias_gen$6

.SUBCKT vias_gen$18
.ENDS vias_gen$18

.SUBCKT nfet$2
.ENDS nfet$2

.SUBCKT vias_gen$7
.ENDS vias_gen$7

.SUBCKT vias_gen$10$1
.ENDS vias_gen$10$1

.SUBCKT vias_gen$2$1$1
.ENDS vias_gen$2$1$1

.SUBCKT pfet$2$1
.ENDS pfet$2$1

.SUBCKT vias_gen$6$1
.ENDS vias_gen$6$1

.SUBCKT vias_gen$18$1
.ENDS vias_gen$18$1

.SUBCKT nfet$2$1
.ENDS nfet$2$1

.SUBCKT vias_gen$7$1
.ENDS vias_gen$7$1

.SUBCKT vias_gen$10$2$1$1$1$1
.ENDS vias_gen$10$2$1$1$1$1

.SUBCKT vias_gen$2$1$2$1$1$1$1
.ENDS vias_gen$2$1$2$1$1$1$1

.SUBCKT pfet$2$2$1$1$1$1
.ENDS pfet$2$2$1$1$1$1

.SUBCKT vias_gen$6$2$1$1$1$1
.ENDS vias_gen$6$2$1$1$1$1

.SUBCKT vias_gen$18$2$1$1$1$1
.ENDS vias_gen$18$2$1$1$1$1

.SUBCKT nfet$2$2$1$1$1$1
.ENDS nfet$2$2$1$1$1$1

.SUBCKT vias_gen$7$2$1$1$1$1
.ENDS vias_gen$7$2$1$1$1$1

.SUBCKT vias_gen$10$1$1$1$1$1$1
.ENDS vias_gen$10$1$1$1$1$1$1

.SUBCKT vias_gen$2$1$1$1$1$1$1$1
.ENDS vias_gen$2$1$1$1$1$1$1$1

.SUBCKT pfet$2$1$1$1$1$1$1
.ENDS pfet$2$1$1$1$1$1$1

.SUBCKT vias_gen$6$1$1$1$1$1$1
.ENDS vias_gen$6$1$1$1$1$1$1

.SUBCKT vias_gen$18$1$1$1$1$1$1
.ENDS vias_gen$18$1$1$1$1$1$1

.SUBCKT nfet$2$1$1$1$1$1$1
.ENDS nfet$2$1$1$1$1$1$1

.SUBCKT vias_gen$7$1$1$1$1$1$1
.ENDS vias_gen$7$1$1$1$1$1$1

.SUBCKT RO_LVT_13St_x1
X$1 RO vias_gen
X$2 RO vias_gen
X$3 RON vias_gen
X$4 RON vias_gen
X$5 RON vias_gen
X$6 RON vias_gen
X$7 RON vias_gen
X$8 GND vias_gen$3
X$9 GND \$36 \$35 VDD sky130_gnd rovcel2_LVT$3$1$1$1$1$1
X$10 GND \$35 \$25 VDD sky130_gnd rovcel2_LVT$2$1$1$1$1$1$1
X$11 GND \$37 \$36 VDD sky130_gnd rovcel2_LVT$2$2$1$1$1$1
X$12 GND \$38 \$37 VDD sky130_gnd rovcel2_LVT$2$1$2$1$1$1
X$13 GND \$39 \$38 VDD sky130_gnd rovcel2_LVT$3$2$1$1$1
X$14 GND \$40 \$39 VDD sky130_gnd rovcel2_LVT$2$1$1$1$2$1
X$15 GND \$41 \$40 VDD sky130_gnd rovcel2_LVT$3$1$1$2$1
X$16 GND \$42 \$41 VDD sky130_gnd rovcel2_LVT$2$2$1$2$1
X$17 GND \$43 \$42 VDD sky130_gnd rovcel2_LVT$2$1$2$2$1
X$18 GND \$44 \$43 VDD sky130_gnd rovcel2_LVT$3$2$2$1
X$19 GND \$45 \$44 VDD sky130_gnd rovcel2_LVT$2$1$1$1$1$2
X$20 GND \$46 \$45 VDD sky130_gnd rovcel2_LVT$3$1$1$1$2
X$21 GND \$47 \$46 VDD sky130_gnd rovcel2_LVT$2$2$1$1$2
X$22 GND \$48 \$47 VDD sky130_gnd rovcel2_LVT$2$1$2$1$2
X$23 GND \$49 \$48 VDD sky130_gnd rovcel2_LVT$3$2$1$2
X$24 GND \$50 \$49 VDD sky130_gnd rovcel2_LVT$2$1$1$1$3
X$25 GND \$51 \$50 VDD sky130_gnd rovcel2_LVT$3$1$1$3
X$26 GND \$52 \$51 VDD sky130_gnd rovcel2_LVT$2$1$1$1$1$1
X$27 GND \$53 \$52 VDD sky130_gnd rovcel2_LVT$3$1$1$1$1
X$28 GND \$54 \$53 VDD sky130_gnd rovcel2_LVT$2$2$1$1$1
X$29 GND \$55 \$54 VDD sky130_gnd rovcel2_LVT$2$1$2$1$1
X$30 GND \$56 \$55 VDD sky130_gnd rovcel2_LVT$3$2$1$1
X$31 GND \$57 \$56 VDD sky130_gnd rovcel2_LVT$2$1$1$1$2
X$32 GND \$58 \$57 VDD sky130_gnd rovcel2_LVT$3$1$1$2
X$33 GND \$59 \$58 VDD sky130_gnd rovcel2_LVT$2$2$1$2
X$34 GND \$60 \$59 VDD sky130_gnd rovcel2_LVT$2$1$2$2
X$35 GND \$61 \$60 VDD sky130_gnd rovcel2_LVT$3$2$2
X$36 GND \$62 \$61 VDD sky130_gnd rovcel2_LVT$2$1$1$1$1
X$37 GND \$63 \$62 VDD sky130_gnd rovcel2_LVT$3$1$1$1
X$38 GND \$64 \$63 VDD sky130_gnd rovcel2_LVT$2$2$1$1
X$39 GND \$65 \$64 VDD sky130_gnd rovcel2_LVT$2$1$2$1
X$40 GND \$66 \$65 VDD sky130_gnd rovcel2_LVT$3$2$1
X$41 GND \$67 \$66 VDD sky130_gnd rovcel2_LVT$2$1$1$1
X$42 GND \$68 \$67 VDD sky130_gnd rovcel2_LVT$3$1$1
X$43 GND \$69 \$68 VDD sky130_gnd rovcel2_LVT$2$2$1
X$44 GND \$70 \$69 VDD sky130_gnd rovcel2_LVT$2$1$2
X$45 GND \$71 \$70 VDD sky130_gnd rovcel2_LVT$3$2
X$46 GND \$72 \$71 VDD sky130_gnd rovcel2_LVT$2$1$1
X$47 GND \$73 \$72 VDD sky130_gnd rovcel2_LVT$3$1
X$48 GND \$74 \$73 VDD sky130_gnd rovcel2_LVT$2$2
X$49 GND \$75 \$74 VDD sky130_gnd rovcel2_LVT$2$1
X$50 GND \$76 \$75 VDD sky130_gnd rovcel2_LVT$3
X$51 GND \$77 \$76 VDD sky130_gnd rovcel2_LVT$2
X$52 GND \$77 VDD sky130_gnd rovcel2_LVT
X$53 GND \$25 \$159 VDD sky130_gnd rovcel2_LVT$1$1$1$1$1$1$1$1
X$54 VDD vias_gen$3
X$55 VDD vias_gen$2
X$56 VDD vias_gen$3
X$57 VDD vias_gen$3
X$58 VDD vias_gen$3
X$59 GND \$159 \$160 VDD sky130_gnd rovcel2_LVT$1$2$1$1$1$1$1
X$60 GND \$160 \$161 VDD sky130_gnd rovcel2_LVT$1$1$2$1$1$1$1
X$61 GND \$161 \$162 VDD sky130_gnd rovcel2_LVT$1$1$1$2$1$1$1
X$62 GND \$162 \$163 VDD sky130_gnd rovcel2_LVT$1$2$2$1$1$1
X$63 GND \$163 \$164 VDD sky130_gnd rovcel2_LVT$1$1$1$1$1$2$1
X$64 GND \$164 \$165 VDD sky130_gnd rovcel2_LVT$1$2$1$1$2$1
X$65 GND \$165 \$166 VDD sky130_gnd rovcel2_LVT$1$1$2$1$2$1
X$66 GND \$166 \$167 VDD sky130_gnd rovcel2_LVT$1$1$1$2$2$1
X$67 GND \$167 \$168 VDD sky130_gnd rovcel2_LVT$1$2$2$2$1
X$68 GND \$168 \$169 VDD sky130_gnd rovcel2_LVT$1$1$1$1$1$1$2
X$69 GND \$169 \$170 VDD sky130_gnd rovcel2_LVT$1$2$1$1$1$2
X$70 GND \$170 \$171 VDD sky130_gnd rovcel2_LVT$1$1$2$1$1$2
X$71 GND \$171 \$172 VDD sky130_gnd rovcel2_LVT$1$1$1$2$1$2
X$72 GND \$172 \$173 VDD sky130_gnd rovcel2_LVT$1$2$2$1$2
X$73 GND \$173 \$174 VDD sky130_gnd rovcel2_LVT$1$1$1$1$1$3
X$74 GND \$174 \$175 VDD sky130_gnd rovcel2_LVT$1$2$1$1$3
X$75 GND \$175 \$176 VDD sky130_gnd rovcel2_LVT$1$1$1$1$1$1$1
X$76 GND \$176 \$177 VDD sky130_gnd rovcel2_LVT$1$2$1$1$1$1
X$77 GND \$177 \$178 VDD sky130_gnd rovcel2_LVT$1$1$2$1$1$1
X$78 GND \$178 \$179 VDD sky130_gnd rovcel2_LVT$1$1$1$2$1$1
X$79 GND \$179 \$180 VDD sky130_gnd rovcel2_LVT$1$2$2$1$1
X$80 GND \$180 \$181 VDD sky130_gnd rovcel2_LVT$1$1$1$1$1$2
X$81 GND \$181 \$182 VDD sky130_gnd rovcel2_LVT$1$2$1$1$2
X$82 GND \$182 \$183 VDD sky130_gnd rovcel2_LVT$1$1$2$1$2
X$83 GND \$183 \$184 VDD sky130_gnd rovcel2_LVT$1$1$1$2$2
X$84 GND \$184 \$185 VDD sky130_gnd rovcel2_LVT$1$2$2$2
X$85 GND \$185 \$186 VDD sky130_gnd rovcel2_LVT$1$1$1$1$1$1
X$86 GND \$186 \$187 VDD sky130_gnd rovcel2_LVT$1$2$1$1$1
X$87 GND \$187 \$188 VDD sky130_gnd rovcel2_LVT$1$1$2$1$1
X$88 GND \$188 \$189 VDD sky130_gnd rovcel2_LVT$1$1$1$2$1
X$89 GND \$189 \$190 VDD sky130_gnd rovcel2_LVT$1$2$2$1
X$90 GND \$190 \$191 VDD sky130_gnd rovcel2_LVT$1$1$1$1$1
X$91 GND \$191 \$192 VDD sky130_gnd rovcel2_LVT$1$2$1$1
X$92 GND \$192 \$193 VDD sky130_gnd rovcel2_LVT$1$1$2$1
X$93 GND \$193 \$194 VDD sky130_gnd rovcel2_LVT$1$1$1$2
X$94 GND \$194 \$195 VDD sky130_gnd rovcel2_LVT$1$2$2
X$95 GND \$195 \$196 VDD sky130_gnd rovcel2_LVT$1$1$1$1
X$96 GND \$196 \$197 VDD sky130_gnd rovcel2_LVT$1$2$1
X$97 GND \$197 \$198 VDD sky130_gnd rovcel2_LVT$1$1$2
X$98 GND \$198 \$199 VDD sky130_gnd rovcel2_LVT$1$1$1
X$99 GND \$199 \$200 VDD sky130_gnd rovcel2_LVT$1$2
X$100 GND \$200 \$201 VDD sky130_gnd rovcel2_LVT$1$1
X$101 GND \$201 \$119 VDD sky130_gnd rovcel2_LVT$1
X$102 GND vias_gen$3
X$103 GND vias_gen$2
M$1 \$78 \$21 \$26 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$2 \$26 \$21 \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$3 \$78 \$21 \$26 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$4 \$26 \$21 \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$5 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$6 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$7 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$8 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$9 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$10 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$11 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$12 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$13 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$14 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$15 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$16 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$17 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$18 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$19 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$20 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$21 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$22 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$23 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$24 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$25 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$26 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$27 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$28 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$29 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$30 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$31 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$32 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$33 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$34 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$35 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$36 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$37 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$38 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$39 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$40 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$41 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$42 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$43 VDD RON \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$44 \$78 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$45 \$80 \$26 \$11 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$46 \$11 \$26 \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$47 \$80 \$26 \$11 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$48 \$11 \$26 \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$49 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$50 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$51 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$52 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$53 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$54 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$55 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$56 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$57 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$58 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$59 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$60 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$61 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$62 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$63 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$64 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$65 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$66 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$67 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$68 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$69 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$70 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$71 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$72 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$73 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$74 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$75 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$76 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$77 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$78 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$79 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$80 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$81 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$82 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$83 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$84 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$85 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$86 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$87 VDD DUT_Footer \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=0.7125 PS=5.05 PD=5.05
M$88 \$80 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=1.425 PS=5.05 PD=10.1
M$89 \$11 RO Drain_Sense VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$90 Drain_Sense RO \$11 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=1.425 PS=5.05 PD=10.1
M$91 \$11 RO Drain_Sense VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$92 Drain_Sense RO \$11 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=1.425 PS=5.05 PD=10.1
M$93 \$11 RO Drain\x20Force VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=1.425 AD=0.7125 PS=10.1 PD=5.05
M$94 Drain\x20Force RO \$11 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=1.425 PS=5.05 PD=10.1
M$95 \$11 RO Drain\x20Force VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=1.425 AD=0.7125 PS=10.1 PD=5.05
M$96 Drain\x20Force RO \$11 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75
+ AS=0.7125 AD=1.425 PS=5.05 PD=10.1
M$97 \$82 \$11 \$27 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$98 \$27 \$11 \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$99 \$82 \$11 \$27 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$100 \$27 \$11 \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$101 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$102 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$103 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$104 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$105 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$106 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$107 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$108 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$109 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$110 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$111 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$112 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$113 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$114 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$115 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$116 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$117 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$118 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$119 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$120 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$121 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$122 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$123 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$124 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$125 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$126 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$127 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$128 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$129 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$130 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$131 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$132 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$133 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$134 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$135 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$136 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$137 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$138 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$139 VDD RON \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=0.7125 PS=5.05 PD=5.05
M$140 \$82 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$141 \$129 VDD \$119 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$142 \$130 VDD \$119 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$143 VDD \$120 \$119 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$144 \$119 \$120 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$145 VDD \$120 \$119 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$146 \$119 \$120 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$147 \$131 VDD \$120 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$148 \$132 VDD \$120 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$149 VDD \$121 \$120 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$150 \$120 \$121 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$151 VDD \$121 \$120 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$152 \$120 \$121 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$153 \$133 VDD \$121 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$154 \$134 VDD \$121 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$155 VDD \$122 \$121 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$156 \$121 \$122 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$157 VDD \$122 \$121 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$158 \$121 \$122 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$159 \$26 RO DUT_Gate VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$160 \$135 VDD \$122 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$161 \$26 RO \$19 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$162 \$136 VDD \$122 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$163 VDD \$123 \$122 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$164 \$122 \$123 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$165 VDD \$123 \$122 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$166 \$122 \$123 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$167 \$137 VDD \$123 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$168 \$138 VDD \$123 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$169 VDD \$124 \$123 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$170 \$123 \$124 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$171 VDD \$124 \$123 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$172 \$123 \$124 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$173 \$139 VDD \$124 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$174 \$140 VDD \$124 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$175 VDD \$125 \$124 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$176 \$124 \$125 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$177 VDD \$125 \$124 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$178 \$124 \$125 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$179 \$141 VDD \$125 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$180 \$142 VDD \$125 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$181 VDD \$126 \$125 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$182 \$125 \$126 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$183 VDD \$126 \$125 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$184 \$125 \$126 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$185 \$143 VDD \$126 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$186 \$144 VDD \$126 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$187 VDD \$127 \$126 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$188 \$126 \$127 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$189 VDD \$127 \$126 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$190 \$126 \$127 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$191 \$145 VDD \$127 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$192 \$146 VDD \$127 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$193 VDD Out \$127 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$194 \$127 Out VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$195 VDD Out \$127 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$196 \$127 Out VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$197 \$147 VDD Out VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$198 \$148 VDD Out VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$199 VDD \$27 Out VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$200 Out \$27 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$201 VDD \$27 Out VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425
+ AD=0.7125 PS=10.1 PD=5.05
M$202 Out \$27 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125
+ AD=1.425 PS=5.05 PD=10.1
M$203 \$27 VDD GND VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$204 \$27 VDD \$20 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
M$205 \$26 \$21 \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$206 \$6 \$21 \$26 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$207 \$6 RO GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$208 GND RO \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$209 \$6 RO GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$210 GND RO \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$211 \$6 RO GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$212 GND RO \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$213 \$6 RO GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$214 GND RO \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$215 \$6 RO GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$216 GND RO \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$217 \$6 RO GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$218 GND RO \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$219 \$6 RO GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$220 GND RO \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$221 \$6 RO GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$222 GND RO \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$223 \$6 RO GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$224 GND RO \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$225 \$6 RO GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$226 GND RO \$6 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$227 \$11 \$26 \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$228 \$12 \$26 \$11 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$229 \$12 DUT_Header GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$230 GND DUT_Header \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$231 \$12 DUT_Header GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$232 GND DUT_Header \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$233 \$12 DUT_Header GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$234 GND DUT_Header \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$235 \$12 DUT_Header GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$236 GND DUT_Header \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$237 \$12 DUT_Header GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$238 GND DUT_Header \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$239 \$12 DUT_Header GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$240 GND DUT_Header \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$241 \$12 DUT_Header GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$242 GND DUT_Header \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$243 \$12 DUT_Header GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$244 GND DUT_Header \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$245 \$12 DUT_Header GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$246 GND DUT_Header \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$247 \$12 DUT_Header GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$248 GND DUT_Header \$12 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$249 \$11 RON Drain_Sense sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$250 Drain_Sense RON \$11 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$251 \$11 RON Drain\x20Force sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35
+ W=2.1 AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$252 Drain\x20Force RON \$11 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35
+ W=2.1 AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$253 \$27 \$11 GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$254 GND \$11 \$27 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$255 \$129 GND \$119 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$256 \$130 GND \$119 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$257 \$119 \$120 GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$258 GND \$120 \$119 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$259 \$131 GND \$120 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$260 \$132 GND \$120 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$261 \$120 \$121 GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$262 GND \$121 \$120 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$263 \$133 GND \$121 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$264 \$134 GND \$121 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$265 \$121 \$122 GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$266 GND \$122 \$121 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$267 \$26 RON DUT_Gate sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$268 \$135 GND \$122 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$269 \$26 RON \$19 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$270 \$136 GND \$122 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$271 \$122 \$123 GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$272 GND \$123 \$122 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$273 \$137 GND \$123 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$274 \$138 GND \$123 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$275 \$123 \$124 GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$276 GND \$124 \$123 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$277 \$139 GND \$124 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$278 \$140 GND \$124 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$279 \$124 \$125 GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$280 GND \$125 \$124 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$281 \$141 GND \$125 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$282 \$142 GND \$125 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$283 \$125 \$126 GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$284 GND \$126 \$125 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$285 \$143 GND \$126 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$286 \$144 GND \$126 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$287 \$126 \$127 GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$288 GND \$127 \$126 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1
+ AS=0.63 AD=0.63 PS=4.8 PD=4.8
M$289 \$145 GND \$127 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$290 \$146 GND \$127 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$291 \$127 Out GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$292 GND Out \$127 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$293 \$147 GND Out sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$294 \$148 GND Out sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$295 Out \$27 GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$296 GND \$27 Out sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$297 \$27 RON GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
M$298 \$27 RON \$20 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45
+ AS=0.135 AD=0.135 PS=1.5 PD=1.5
.ENDS RO_LVT_13St_x1

.SUBCKT rovcel2_LVT$2$1$1$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$1$1$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$1$1$1$1$1
X$3 IN OUT GND nfet$5$1$1$1$1$1$1
X$4 IN GND OUT nfet$5$1$1$1$1$1$1
X$5 GND vias_gen$17$2$1$1$1$1$1$1
X$6 GND vias_gen$17$2$1$1$1$1$1$1
X$7 GND vias_gen$15$2$1$1$1$1$1$1
X$8 OUT vias_gen$12$2$1$1$1$1$1$1
X$9 OUT vias_gen$8$2$1$1$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$2$1$1$1$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$2$1$1$1$1$1$1
X$12 OUT vias_gen$8$2$1$1$1$1$1$1
X$13 OUT vias_gen$12$2$1$1$1$1$1$1
X$14 IN OUT VDD VDD pfet$4$2$1$1$1$1$1$1
X$15 IN VDD OUT VDD pfet$4$2$1$1$1$1$1$1
X$16 OUT vias_gen$13$2$1$1$1$1$1$1
X$17 IN VDD OUT VDD pfet$4$2$1$1$1$1$1$1
X$18 OUT vias_gen$13$2$1$1$1$1$1$1
X$19 IN OUT VDD VDD pfet$4$2$1$1$1$1$1$1
X$20 OUT vias_gen$16$2$1$1$1$1$1$1
X$21 OUT vias_gen$16$2$1$1$1$1$1$1
X$22 IN vias_gen$14$2$1$1$1$1$1$1
X$23 IN vias_gen$14$2$1$1$1$1$1$1
X$24 IN vias_gen$14$2$1$1$1$1$1$1
X$25 IN vias_gen$14$2$1$1$1$1$1$1
X$26 VDD vias_gen$17$2$1$1$1$1$1$1
X$27 VDD vias_gen$17$2$1$1$1$1$1$1
X$28 VDD vias_gen$15$2$1$1$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$1$1$1$1$1

.SUBCKT rovcel2_LVT$1$1$1$1$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$1$1$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$1$1$1$1$1
X$3 IN GND OUT nfet$4$1$1$1$1$1$1$1
X$4 GND vias_gen$17$1$1$1$1$1$1$1$1
X$5 GND vias_gen$15$1$1$1$1$1$1$1$1
X$6 GND vias_gen$17$1$1$1$1$1$1$1$1
X$7 IN OUT GND nfet$4$1$1$1$1$1$1$1
X$8 OUT vias_gen$12$1$1$1$1$1$1$1$1
X$9 OUT vias_gen$8$1$1$1$1$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$1$1$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$1$1$1$1$1
X$12 OUT vias_gen$8$1$1$1$1$1$1$1$1
X$13 OUT vias_gen$12$1$1$1$1$1$1$1$1
X$14 OUT vias_gen$16$1$1$1$1$1$1$1$1
X$15 OUT vias_gen$16$1$1$1$1$1$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$1$1$1$1$1$1
X$17 OUT vias_gen$13$1$1$1$1$1$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$1$1$1$1$1$1
X$19 OUT vias_gen$13$1$1$1$1$1$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$1$1$1$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$1$1$1$1$1$1
X$22 IN vias_gen$14$1$1$1$1$1$1$1$1
X$23 IN vias_gen$14$1$1$1$1$1$1$1$1
X$24 IN vias_gen$14$1$1$1$1$1$1$1$1
X$25 IN vias_gen$14$1$1$1$1$1$1$1$1
X$26 VDD vias_gen$17$1$1$1$1$1$1$1$1
X$27 VDD vias_gen$15$1$1$1$1$1$1$1$1
X$28 VDD vias_gen$17$1$1$1$1$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$1$1$1$1$1

.SUBCKT rovcel2_LVT$3$1$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$1$1$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$1$1$1$1$1
X$3 IN OUT GND nfet$6$1$1$1$1$1
X$4 IN GND OUT nfet$6$1$1$1$1$1
X$5 GND vias_gen$17$3$1$1$1$1$1
X$6 GND vias_gen$17$3$1$1$1$1$1
X$7 GND vias_gen$15$3$1$1$1$1$1
X$8 OUT vias_gen$12$3$1$1$1$1$1
X$9 OUT vias_gen$8$3$1$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$3$1$1$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$3$1$1$1$1$1
X$12 OUT vias_gen$8$3$1$1$1$1$1
X$13 OUT vias_gen$12$3$1$1$1$1$1
X$14 IN OUT VDD VDD pfet$4$3$1$1$1$1$1
X$15 IN VDD OUT VDD pfet$4$3$1$1$1$1$1
X$16 OUT vias_gen$13$3$1$1$1$1$1
X$17 IN VDD OUT VDD pfet$4$3$1$1$1$1$1
X$18 OUT vias_gen$13$3$1$1$1$1$1
X$19 IN OUT VDD VDD pfet$4$3$1$1$1$1$1
X$20 OUT vias_gen$16$3$1$1$1$1$1
X$21 OUT vias_gen$16$3$1$1$1$1$1
X$22 IN vias_gen$14$3$1$1$1$1$1
X$23 IN vias_gen$14$3$1$1$1$1$1
X$24 IN vias_gen$14$3$1$1$1$1$1
X$25 IN vias_gen$14$3$1$1$1$1$1
X$26 VDD vias_gen$17$3$1$1$1$1$1
X$27 VDD vias_gen$17$3$1$1$1$1$1
X$28 VDD vias_gen$15$3$1$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$1$1$1$1$1

.SUBCKT rovcel2_LVT$1$2$1$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$1$1$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$1$1$1$1$1
X$3 IN GND OUT nfet$4$2$1$1$1$1$1
X$4 GND vias_gen$17$1$2$1$1$1$1$1
X$5 GND vias_gen$15$1$2$1$1$1$1$1
X$6 GND vias_gen$17$1$2$1$1$1$1$1
X$7 IN OUT GND nfet$4$2$1$1$1$1$1
X$8 OUT vias_gen$12$1$2$1$1$1$1$1
X$9 OUT vias_gen$8$1$2$1$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$2$1$1$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$2$1$1$1$1$1
X$12 OUT vias_gen$8$1$2$1$1$1$1$1
X$13 OUT vias_gen$12$1$2$1$1$1$1$1
X$14 OUT vias_gen$16$1$2$1$1$1$1$1
X$15 OUT vias_gen$16$1$2$1$1$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$2$1$1$1$1$1
X$17 OUT vias_gen$13$1$2$1$1$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$2$1$1$1$1$1
X$19 OUT vias_gen$13$1$2$1$1$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$2$1$1$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$2$1$1$1$1$1
X$22 IN vias_gen$14$1$2$1$1$1$1$1
X$23 IN vias_gen$14$1$2$1$1$1$1$1
X$24 IN vias_gen$14$1$2$1$1$1$1$1
X$25 IN vias_gen$14$1$2$1$1$1$1$1
X$26 VDD vias_gen$17$1$2$1$1$1$1$1
X$27 VDD vias_gen$15$1$2$1$1$1$1$1
X$28 VDD vias_gen$17$1$2$1$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$1$1$1$1$1

.SUBCKT rovcel2_LVT$2$2$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$2$1$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$2$1$1$1$1
X$3 IN OUT GND nfet$5$2$1$1$1$1
X$4 IN GND OUT nfet$5$2$1$1$1$1
X$5 GND vias_gen$17$2$2$1$1$1$1
X$6 GND vias_gen$17$2$2$1$1$1$1
X$7 GND vias_gen$15$2$2$1$1$1$1
X$8 OUT vias_gen$12$2$2$1$1$1$1
X$9 OUT vias_gen$8$2$2$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$2$2$1$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$2$2$1$1$1$1
X$12 OUT vias_gen$8$2$2$1$1$1$1
X$13 OUT vias_gen$12$2$2$1$1$1$1
X$14 IN OUT VDD VDD pfet$4$2$2$1$1$1$1
X$15 IN VDD OUT VDD pfet$4$2$2$1$1$1$1
X$16 OUT vias_gen$13$2$2$1$1$1$1
X$17 IN VDD OUT VDD pfet$4$2$2$1$1$1$1
X$18 OUT vias_gen$13$2$2$1$1$1$1
X$19 IN OUT VDD VDD pfet$4$2$2$1$1$1$1
X$20 OUT vias_gen$16$2$2$1$1$1$1
X$21 OUT vias_gen$16$2$2$1$1$1$1
X$22 IN vias_gen$14$2$2$1$1$1$1
X$23 IN vias_gen$14$2$2$1$1$1$1
X$24 IN vias_gen$14$2$2$1$1$1$1
X$25 IN vias_gen$14$2$2$1$1$1$1
X$26 VDD vias_gen$17$2$2$1$1$1$1
X$27 VDD vias_gen$17$2$2$1$1$1$1
X$28 VDD vias_gen$15$2$2$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$2$1$1$1$1

.SUBCKT rovcel2_LVT$1$1$2$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$2$1$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$2$1$1$1$1
X$3 IN GND OUT nfet$4$1$2$1$1$1$1
X$4 GND vias_gen$17$1$1$2$1$1$1$1
X$5 GND vias_gen$15$1$1$2$1$1$1$1
X$6 GND vias_gen$17$1$1$2$1$1$1$1
X$7 IN OUT GND nfet$4$1$2$1$1$1$1
X$8 OUT vias_gen$12$1$1$2$1$1$1$1
X$9 OUT vias_gen$8$1$1$2$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$2$1$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$2$1$1$1$1
X$12 OUT vias_gen$8$1$1$2$1$1$1$1
X$13 OUT vias_gen$12$1$1$2$1$1$1$1
X$14 OUT vias_gen$16$1$1$2$1$1$1$1
X$15 OUT vias_gen$16$1$1$2$1$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$2$1$1$1$1
X$17 OUT vias_gen$13$1$1$2$1$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$2$1$1$1$1
X$19 OUT vias_gen$13$1$1$2$1$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$2$1$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$2$1$1$1$1
X$22 IN vias_gen$14$1$1$2$1$1$1$1
X$23 IN vias_gen$14$1$1$2$1$1$1$1
X$24 IN vias_gen$14$1$1$2$1$1$1$1
X$25 IN vias_gen$14$1$1$2$1$1$1$1
X$26 VDD vias_gen$17$1$1$2$1$1$1$1
X$27 VDD vias_gen$15$1$1$2$1$1$1$1
X$28 VDD vias_gen$17$1$1$2$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$2$1$1$1$1

.SUBCKT rovcel2_LVT$2$1$2$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$2$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$2$1$1$1
X$3 IN OUT GND nfet$5$1$2$1$1$1
X$4 IN GND OUT nfet$5$1$2$1$1$1
X$5 GND vias_gen$17$2$1$2$1$1$1
X$6 GND vias_gen$17$2$1$2$1$1$1
X$7 GND vias_gen$15$2$1$2$1$1$1
X$8 OUT vias_gen$12$2$1$2$1$1$1
X$9 OUT vias_gen$8$2$1$2$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$2$1$2$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$2$1$2$1$1$1
X$12 OUT vias_gen$8$2$1$2$1$1$1
X$13 OUT vias_gen$12$2$1$2$1$1$1
X$14 IN OUT VDD VDD pfet$4$2$1$2$1$1$1
X$15 IN VDD OUT VDD pfet$4$2$1$2$1$1$1
X$16 OUT vias_gen$13$2$1$2$1$1$1
X$17 IN VDD OUT VDD pfet$4$2$1$2$1$1$1
X$18 OUT vias_gen$13$2$1$2$1$1$1
X$19 IN OUT VDD VDD pfet$4$2$1$2$1$1$1
X$20 OUT vias_gen$16$2$1$2$1$1$1
X$21 OUT vias_gen$16$2$1$2$1$1$1
X$22 IN vias_gen$14$2$1$2$1$1$1
X$23 IN vias_gen$14$2$1$2$1$1$1
X$24 IN vias_gen$14$2$1$2$1$1$1
X$25 IN vias_gen$14$2$1$2$1$1$1
X$26 VDD vias_gen$17$2$1$2$1$1$1
X$27 VDD vias_gen$17$2$1$2$1$1$1
X$28 VDD vias_gen$15$2$1$2$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$2$1$1$1

.SUBCKT rovcel2_LVT$1$1$1$2$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$2$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$2$1$1$1
X$3 IN GND OUT nfet$4$1$1$2$1$1$1
X$4 GND vias_gen$17$1$1$1$2$1$1$1
X$5 GND vias_gen$15$1$1$1$2$1$1$1
X$6 GND vias_gen$17$1$1$1$2$1$1$1
X$7 IN OUT GND nfet$4$1$1$2$1$1$1
X$8 OUT vias_gen$12$1$1$1$2$1$1$1
X$9 OUT vias_gen$8$1$1$1$2$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$2$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$2$1$1$1
X$12 OUT vias_gen$8$1$1$1$2$1$1$1
X$13 OUT vias_gen$12$1$1$1$2$1$1$1
X$14 OUT vias_gen$16$1$1$1$2$1$1$1
X$15 OUT vias_gen$16$1$1$1$2$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$1$2$1$1$1
X$17 OUT vias_gen$13$1$1$1$2$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$1$2$1$1$1
X$19 OUT vias_gen$13$1$1$1$2$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$1$2$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$1$2$1$1$1
X$22 IN vias_gen$14$1$1$1$2$1$1$1
X$23 IN vias_gen$14$1$1$1$2$1$1$1
X$24 IN vias_gen$14$1$1$1$2$1$1$1
X$25 IN vias_gen$14$1$1$1$2$1$1$1
X$26 VDD vias_gen$17$1$1$1$2$1$1$1
X$27 VDD vias_gen$15$1$1$1$2$1$1$1
X$28 VDD vias_gen$17$1$1$1$2$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$2$1$1$1

.SUBCKT rovcel2_LVT$3$2$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$2$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$2$1$1$1
X$3 IN OUT GND nfet$6$2$1$1$1
X$4 IN GND OUT nfet$6$2$1$1$1
X$5 GND vias_gen$17$3$2$1$1$1
X$6 GND vias_gen$17$3$2$1$1$1
X$7 GND vias_gen$15$3$2$1$1$1
X$8 OUT vias_gen$12$3$2$1$1$1
X$9 OUT vias_gen$8$3$2$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$3$2$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$3$2$1$1$1
X$12 OUT vias_gen$8$3$2$1$1$1
X$13 OUT vias_gen$12$3$2$1$1$1
X$14 IN OUT VDD VDD pfet$4$3$2$1$1$1
X$15 IN VDD OUT VDD pfet$4$3$2$1$1$1
X$16 OUT vias_gen$13$3$2$1$1$1
X$17 IN VDD OUT VDD pfet$4$3$2$1$1$1
X$18 OUT vias_gen$13$3$2$1$1$1
X$19 IN OUT VDD VDD pfet$4$3$2$1$1$1
X$20 OUT vias_gen$16$3$2$1$1$1
X$21 OUT vias_gen$16$3$2$1$1$1
X$22 IN vias_gen$14$3$2$1$1$1
X$23 IN vias_gen$14$3$2$1$1$1
X$24 IN vias_gen$14$3$2$1$1$1
X$25 IN vias_gen$14$3$2$1$1$1
X$26 VDD vias_gen$17$3$2$1$1$1
X$27 VDD vias_gen$17$3$2$1$1$1
X$28 VDD vias_gen$15$3$2$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$2$1$1$1

.SUBCKT rovcel2_LVT$1$2$2$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$2$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$2$1$1$1
X$3 IN GND OUT nfet$4$2$2$1$1$1
X$4 GND vias_gen$17$1$2$2$1$1$1
X$5 GND vias_gen$15$1$2$2$1$1$1
X$6 GND vias_gen$17$1$2$2$1$1$1
X$7 IN OUT GND nfet$4$2$2$1$1$1
X$8 OUT vias_gen$12$1$2$2$1$1$1
X$9 OUT vias_gen$8$1$2$2$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$2$2$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$2$2$1$1$1
X$12 OUT vias_gen$8$1$2$2$1$1$1
X$13 OUT vias_gen$12$1$2$2$1$1$1
X$14 OUT vias_gen$16$1$2$2$1$1$1
X$15 OUT vias_gen$16$1$2$2$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$2$2$1$1$1
X$17 OUT vias_gen$13$1$2$2$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$2$2$1$1$1
X$19 OUT vias_gen$13$1$2$2$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$2$2$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$2$2$1$1$1
X$22 IN vias_gen$14$1$2$2$1$1$1
X$23 IN vias_gen$14$1$2$2$1$1$1
X$24 IN vias_gen$14$1$2$2$1$1$1
X$25 IN vias_gen$14$1$2$2$1$1$1
X$26 VDD vias_gen$17$1$2$2$1$1$1
X$27 VDD vias_gen$15$1$2$2$1$1$1
X$28 VDD vias_gen$17$1$2$2$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$2$1$1$1

.SUBCKT rovcel2_LVT$2$1$1$1$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$1$1$2$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$1$1$2$1
X$3 IN OUT GND nfet$5$1$1$1$2$1
X$4 IN GND OUT nfet$5$1$1$1$2$1
X$5 GND vias_gen$17$2$1$1$1$2$1
X$6 GND vias_gen$17$2$1$1$1$2$1
X$7 GND vias_gen$15$2$1$1$1$2$1
X$8 OUT vias_gen$12$2$1$1$1$2$1
X$9 OUT vias_gen$8$2$1$1$1$2$1
X$10 VDD VDD \$25 OUT pfet$5$2$1$1$1$2$1
X$11 VDD VDD \$28 OUT pfet$5$2$1$1$1$2$1
X$12 OUT vias_gen$8$2$1$1$1$2$1
X$13 OUT vias_gen$12$2$1$1$1$2$1
X$14 IN OUT VDD VDD pfet$4$2$1$1$1$2$1
X$15 IN VDD OUT VDD pfet$4$2$1$1$1$2$1
X$16 OUT vias_gen$13$2$1$1$1$2$1
X$17 IN VDD OUT VDD pfet$4$2$1$1$1$2$1
X$18 OUT vias_gen$13$2$1$1$1$2$1
X$19 IN OUT VDD VDD pfet$4$2$1$1$1$2$1
X$20 OUT vias_gen$16$2$1$1$1$2$1
X$21 OUT vias_gen$16$2$1$1$1$2$1
X$22 IN vias_gen$14$2$1$1$1$2$1
X$23 IN vias_gen$14$2$1$1$1$2$1
X$24 IN vias_gen$14$2$1$1$1$2$1
X$25 IN vias_gen$14$2$1$1$1$2$1
X$26 VDD vias_gen$17$2$1$1$1$2$1
X$27 VDD vias_gen$17$2$1$1$1$2$1
X$28 VDD vias_gen$15$2$1$1$1$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$1$1$2$1

.SUBCKT rovcel2_LVT$1$1$1$1$1$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$1$1$2$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$1$1$2$1
X$3 IN GND OUT nfet$4$1$1$1$1$2$1
X$4 GND vias_gen$17$1$1$1$1$1$2$1
X$5 GND vias_gen$15$1$1$1$1$1$2$1
X$6 GND vias_gen$17$1$1$1$1$1$2$1
X$7 IN OUT GND nfet$4$1$1$1$1$2$1
X$8 OUT vias_gen$12$1$1$1$1$1$2$1
X$9 OUT vias_gen$8$1$1$1$1$1$2$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$1$1$2$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$1$1$2$1
X$12 OUT vias_gen$8$1$1$1$1$1$2$1
X$13 OUT vias_gen$12$1$1$1$1$1$2$1
X$14 OUT vias_gen$16$1$1$1$1$1$2$1
X$15 OUT vias_gen$16$1$1$1$1$1$2$1
X$16 IN OUT VDD VDD pfet$4$1$1$1$1$1$2$1
X$17 OUT vias_gen$13$1$1$1$1$1$2$1
X$18 IN VDD OUT VDD pfet$4$1$1$1$1$1$2$1
X$19 OUT vias_gen$13$1$1$1$1$1$2$1
X$20 IN VDD OUT VDD pfet$4$1$1$1$1$1$2$1
X$21 IN OUT VDD VDD pfet$4$1$1$1$1$1$2$1
X$22 IN vias_gen$14$1$1$1$1$1$2$1
X$23 IN vias_gen$14$1$1$1$1$1$2$1
X$24 IN vias_gen$14$1$1$1$1$1$2$1
X$25 IN vias_gen$14$1$1$1$1$1$2$1
X$26 VDD vias_gen$17$1$1$1$1$1$2$1
X$27 VDD vias_gen$15$1$1$1$1$1$2$1
X$28 VDD vias_gen$17$1$1$1$1$1$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$1$1$2$1

.SUBCKT rovcel2_LVT$3$1$1$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$1$1$2$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$1$1$2$1
X$3 IN OUT GND nfet$6$1$1$2$1
X$4 IN GND OUT nfet$6$1$1$2$1
X$5 GND vias_gen$17$3$1$1$2$1
X$6 GND vias_gen$17$3$1$1$2$1
X$7 GND vias_gen$15$3$1$1$2$1
X$8 OUT vias_gen$12$3$1$1$2$1
X$9 OUT vias_gen$8$3$1$1$2$1
X$10 VDD VDD \$25 OUT pfet$5$3$1$1$2$1
X$11 VDD VDD \$28 OUT pfet$5$3$1$1$2$1
X$12 OUT vias_gen$8$3$1$1$2$1
X$13 OUT vias_gen$12$3$1$1$2$1
X$14 IN OUT VDD VDD pfet$4$3$1$1$2$1
X$15 IN VDD OUT VDD pfet$4$3$1$1$2$1
X$16 OUT vias_gen$13$3$1$1$2$1
X$17 IN VDD OUT VDD pfet$4$3$1$1$2$1
X$18 OUT vias_gen$13$3$1$1$2$1
X$19 IN OUT VDD VDD pfet$4$3$1$1$2$1
X$20 OUT vias_gen$16$3$1$1$2$1
X$21 OUT vias_gen$16$3$1$1$2$1
X$22 IN vias_gen$14$3$1$1$2$1
X$23 IN vias_gen$14$3$1$1$2$1
X$24 IN vias_gen$14$3$1$1$2$1
X$25 IN vias_gen$14$3$1$1$2$1
X$26 VDD vias_gen$17$3$1$1$2$1
X$27 VDD vias_gen$17$3$1$1$2$1
X$28 VDD vias_gen$15$3$1$1$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$1$1$2$1

.SUBCKT rovcel2_LVT$1$2$1$1$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$1$1$2$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$1$1$2$1
X$3 IN GND OUT nfet$4$2$1$1$2$1
X$4 GND vias_gen$17$1$2$1$1$2$1
X$5 GND vias_gen$15$1$2$1$1$2$1
X$6 GND vias_gen$17$1$2$1$1$2$1
X$7 IN OUT GND nfet$4$2$1$1$2$1
X$8 OUT vias_gen$12$1$2$1$1$2$1
X$9 OUT vias_gen$8$1$2$1$1$2$1
X$10 VDD VDD \$25 OUT pfet$5$1$2$1$1$2$1
X$11 VDD VDD \$27 OUT pfet$5$1$2$1$1$2$1
X$12 OUT vias_gen$8$1$2$1$1$2$1
X$13 OUT vias_gen$12$1$2$1$1$2$1
X$14 OUT vias_gen$16$1$2$1$1$2$1
X$15 OUT vias_gen$16$1$2$1$1$2$1
X$16 IN OUT VDD VDD pfet$4$1$2$1$1$2$1
X$17 OUT vias_gen$13$1$2$1$1$2$1
X$18 IN VDD OUT VDD pfet$4$1$2$1$1$2$1
X$19 OUT vias_gen$13$1$2$1$1$2$1
X$20 IN VDD OUT VDD pfet$4$1$2$1$1$2$1
X$21 IN OUT VDD VDD pfet$4$1$2$1$1$2$1
X$22 IN vias_gen$14$1$2$1$1$2$1
X$23 IN vias_gen$14$1$2$1$1$2$1
X$24 IN vias_gen$14$1$2$1$1$2$1
X$25 IN vias_gen$14$1$2$1$1$2$1
X$26 VDD vias_gen$17$1$2$1$1$2$1
X$27 VDD vias_gen$15$1$2$1$1$2$1
X$28 VDD vias_gen$17$1$2$1$1$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$1$1$2$1

.SUBCKT rovcel2_LVT$2$2$1$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$2$1$2$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$2$1$2$1
X$3 IN OUT GND nfet$5$2$1$2$1
X$4 IN GND OUT nfet$5$2$1$2$1
X$5 GND vias_gen$17$2$2$1$2$1
X$6 GND vias_gen$17$2$2$1$2$1
X$7 GND vias_gen$15$2$2$1$2$1
X$8 OUT vias_gen$12$2$2$1$2$1
X$9 OUT vias_gen$8$2$2$1$2$1
X$10 VDD VDD \$25 OUT pfet$5$2$2$1$2$1
X$11 VDD VDD \$28 OUT pfet$5$2$2$1$2$1
X$12 OUT vias_gen$8$2$2$1$2$1
X$13 OUT vias_gen$12$2$2$1$2$1
X$14 IN OUT VDD VDD pfet$4$2$2$1$2$1
X$15 IN VDD OUT VDD pfet$4$2$2$1$2$1
X$16 OUT vias_gen$13$2$2$1$2$1
X$17 IN VDD OUT VDD pfet$4$2$2$1$2$1
X$18 OUT vias_gen$13$2$2$1$2$1
X$19 IN OUT VDD VDD pfet$4$2$2$1$2$1
X$20 OUT vias_gen$16$2$2$1$2$1
X$21 OUT vias_gen$16$2$2$1$2$1
X$22 IN vias_gen$14$2$2$1$2$1
X$23 IN vias_gen$14$2$2$1$2$1
X$24 IN vias_gen$14$2$2$1$2$1
X$25 IN vias_gen$14$2$2$1$2$1
X$26 VDD vias_gen$17$2$2$1$2$1
X$27 VDD vias_gen$17$2$2$1$2$1
X$28 VDD vias_gen$15$2$2$1$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$2$1$2$1

.SUBCKT rovcel2_LVT$1$1$2$1$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$2$1$2$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$2$1$2$1
X$3 IN GND OUT nfet$4$1$2$1$2$1
X$4 GND vias_gen$17$1$1$2$1$2$1
X$5 GND vias_gen$15$1$1$2$1$2$1
X$6 GND vias_gen$17$1$1$2$1$2$1
X$7 IN OUT GND nfet$4$1$2$1$2$1
X$8 OUT vias_gen$12$1$1$2$1$2$1
X$9 OUT vias_gen$8$1$1$2$1$2$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$2$1$2$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$2$1$2$1
X$12 OUT vias_gen$8$1$1$2$1$2$1
X$13 OUT vias_gen$12$1$1$2$1$2$1
X$14 OUT vias_gen$16$1$1$2$1$2$1
X$15 OUT vias_gen$16$1$1$2$1$2$1
X$16 IN OUT VDD VDD pfet$4$1$1$2$1$2$1
X$17 OUT vias_gen$13$1$1$2$1$2$1
X$18 IN VDD OUT VDD pfet$4$1$1$2$1$2$1
X$19 OUT vias_gen$13$1$1$2$1$2$1
X$20 IN VDD OUT VDD pfet$4$1$1$2$1$2$1
X$21 IN OUT VDD VDD pfet$4$1$1$2$1$2$1
X$22 IN vias_gen$14$1$1$2$1$2$1
X$23 IN vias_gen$14$1$1$2$1$2$1
X$24 IN vias_gen$14$1$1$2$1$2$1
X$25 IN vias_gen$14$1$1$2$1$2$1
X$26 VDD vias_gen$17$1$1$2$1$2$1
X$27 VDD vias_gen$15$1$1$2$1$2$1
X$28 VDD vias_gen$17$1$1$2$1$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$2$1$2$1

.SUBCKT rovcel2_LVT$2$1$2$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$2$2$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$2$2$1
X$3 IN OUT GND nfet$5$1$2$2$1
X$4 IN GND OUT nfet$5$1$2$2$1
X$5 GND vias_gen$17$2$1$2$2$1
X$6 GND vias_gen$17$2$1$2$2$1
X$7 GND vias_gen$15$2$1$2$2$1
X$8 OUT vias_gen$12$2$1$2$2$1
X$9 OUT vias_gen$8$2$1$2$2$1
X$10 VDD VDD \$25 OUT pfet$5$2$1$2$2$1
X$11 VDD VDD \$28 OUT pfet$5$2$1$2$2$1
X$12 OUT vias_gen$8$2$1$2$2$1
X$13 OUT vias_gen$12$2$1$2$2$1
X$14 IN OUT VDD VDD pfet$4$2$1$2$2$1
X$15 IN VDD OUT VDD pfet$4$2$1$2$2$1
X$16 OUT vias_gen$13$2$1$2$2$1
X$17 IN VDD OUT VDD pfet$4$2$1$2$2$1
X$18 OUT vias_gen$13$2$1$2$2$1
X$19 IN OUT VDD VDD pfet$4$2$1$2$2$1
X$20 OUT vias_gen$16$2$1$2$2$1
X$21 OUT vias_gen$16$2$1$2$2$1
X$22 IN vias_gen$14$2$1$2$2$1
X$23 IN vias_gen$14$2$1$2$2$1
X$24 IN vias_gen$14$2$1$2$2$1
X$25 IN vias_gen$14$2$1$2$2$1
X$26 VDD vias_gen$17$2$1$2$2$1
X$27 VDD vias_gen$17$2$1$2$2$1
X$28 VDD vias_gen$15$2$1$2$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$2$2$1

.SUBCKT rovcel2_LVT$1$1$1$2$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$2$2$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$2$2$1
X$3 IN GND OUT nfet$4$1$1$2$2$1
X$4 GND vias_gen$17$1$1$1$2$2$1
X$5 GND vias_gen$15$1$1$1$2$2$1
X$6 GND vias_gen$17$1$1$1$2$2$1
X$7 IN OUT GND nfet$4$1$1$2$2$1
X$8 OUT vias_gen$12$1$1$1$2$2$1
X$9 OUT vias_gen$8$1$1$1$2$2$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$2$2$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$2$2$1
X$12 OUT vias_gen$8$1$1$1$2$2$1
X$13 OUT vias_gen$12$1$1$1$2$2$1
X$14 OUT vias_gen$16$1$1$1$2$2$1
X$15 OUT vias_gen$16$1$1$1$2$2$1
X$16 IN OUT VDD VDD pfet$4$1$1$1$2$2$1
X$17 OUT vias_gen$13$1$1$1$2$2$1
X$18 IN VDD OUT VDD pfet$4$1$1$1$2$2$1
X$19 OUT vias_gen$13$1$1$1$2$2$1
X$20 IN VDD OUT VDD pfet$4$1$1$1$2$2$1
X$21 IN OUT VDD VDD pfet$4$1$1$1$2$2$1
X$22 IN vias_gen$14$1$1$1$2$2$1
X$23 IN vias_gen$14$1$1$1$2$2$1
X$24 IN vias_gen$14$1$1$1$2$2$1
X$25 IN vias_gen$14$1$1$1$2$2$1
X$26 VDD vias_gen$17$1$1$1$2$2$1
X$27 VDD vias_gen$15$1$1$1$2$2$1
X$28 VDD vias_gen$17$1$1$1$2$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$2$2$1

.SUBCKT rovcel2_LVT$3$2$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$2$2$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$2$2$1
X$3 IN OUT GND nfet$6$2$2$1
X$4 IN GND OUT nfet$6$2$2$1
X$5 GND vias_gen$17$3$2$2$1
X$6 GND vias_gen$17$3$2$2$1
X$7 GND vias_gen$15$3$2$2$1
X$8 OUT vias_gen$12$3$2$2$1
X$9 OUT vias_gen$8$3$2$2$1
X$10 VDD VDD \$25 OUT pfet$5$3$2$2$1
X$11 VDD VDD \$28 OUT pfet$5$3$2$2$1
X$12 OUT vias_gen$8$3$2$2$1
X$13 OUT vias_gen$12$3$2$2$1
X$14 IN OUT VDD VDD pfet$4$3$2$2$1
X$15 IN VDD OUT VDD pfet$4$3$2$2$1
X$16 OUT vias_gen$13$3$2$2$1
X$17 IN VDD OUT VDD pfet$4$3$2$2$1
X$18 OUT vias_gen$13$3$2$2$1
X$19 IN OUT VDD VDD pfet$4$3$2$2$1
X$20 OUT vias_gen$16$3$2$2$1
X$21 OUT vias_gen$16$3$2$2$1
X$22 IN vias_gen$14$3$2$2$1
X$23 IN vias_gen$14$3$2$2$1
X$24 IN vias_gen$14$3$2$2$1
X$25 IN vias_gen$14$3$2$2$1
X$26 VDD vias_gen$17$3$2$2$1
X$27 VDD vias_gen$17$3$2$2$1
X$28 VDD vias_gen$15$3$2$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$2$2$1

.SUBCKT rovcel2_LVT$1$2$2$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$2$2$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$2$2$1
X$3 IN GND OUT nfet$4$2$2$2$1
X$4 GND vias_gen$17$1$2$2$2$1
X$5 GND vias_gen$15$1$2$2$2$1
X$6 GND vias_gen$17$1$2$2$2$1
X$7 IN OUT GND nfet$4$2$2$2$1
X$8 OUT vias_gen$12$1$2$2$2$1
X$9 OUT vias_gen$8$1$2$2$2$1
X$10 VDD VDD \$25 OUT pfet$5$1$2$2$2$1
X$11 VDD VDD \$27 OUT pfet$5$1$2$2$2$1
X$12 OUT vias_gen$8$1$2$2$2$1
X$13 OUT vias_gen$12$1$2$2$2$1
X$14 OUT vias_gen$16$1$2$2$2$1
X$15 OUT vias_gen$16$1$2$2$2$1
X$16 IN OUT VDD VDD pfet$4$1$2$2$2$1
X$17 OUT vias_gen$13$1$2$2$2$1
X$18 IN VDD OUT VDD pfet$4$1$2$2$2$1
X$19 OUT vias_gen$13$1$2$2$2$1
X$20 IN VDD OUT VDD pfet$4$1$2$2$2$1
X$21 IN OUT VDD VDD pfet$4$1$2$2$2$1
X$22 IN vias_gen$14$1$2$2$2$1
X$23 IN vias_gen$14$1$2$2$2$1
X$24 IN vias_gen$14$1$2$2$2$1
X$25 IN vias_gen$14$1$2$2$2$1
X$26 VDD vias_gen$17$1$2$2$2$1
X$27 VDD vias_gen$15$1$2$2$2$1
X$28 VDD vias_gen$17$1$2$2$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$2$2$1

.SUBCKT rovcel2_LVT$2$1$1$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$1$1$1$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$1$1$1$2
X$3 IN OUT GND nfet$5$1$1$1$1$2
X$4 IN GND OUT nfet$5$1$1$1$1$2
X$5 GND vias_gen$17$2$1$1$1$1$2
X$6 GND vias_gen$17$2$1$1$1$1$2
X$7 GND vias_gen$15$2$1$1$1$1$2
X$8 OUT vias_gen$12$2$1$1$1$1$2
X$9 OUT vias_gen$8$2$1$1$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$2$1$1$1$1$2
X$11 VDD VDD \$28 OUT pfet$5$2$1$1$1$1$2
X$12 OUT vias_gen$8$2$1$1$1$1$2
X$13 OUT vias_gen$12$2$1$1$1$1$2
X$14 IN OUT VDD VDD pfet$4$2$1$1$1$1$2
X$15 IN VDD OUT VDD pfet$4$2$1$1$1$1$2
X$16 OUT vias_gen$13$2$1$1$1$1$2
X$17 IN VDD OUT VDD pfet$4$2$1$1$1$1$2
X$18 OUT vias_gen$13$2$1$1$1$1$2
X$19 IN OUT VDD VDD pfet$4$2$1$1$1$1$2
X$20 OUT vias_gen$16$2$1$1$1$1$2
X$21 OUT vias_gen$16$2$1$1$1$1$2
X$22 IN vias_gen$14$2$1$1$1$1$2
X$23 IN vias_gen$14$2$1$1$1$1$2
X$24 IN vias_gen$14$2$1$1$1$1$2
X$25 IN vias_gen$14$2$1$1$1$1$2
X$26 VDD vias_gen$17$2$1$1$1$1$2
X$27 VDD vias_gen$17$2$1$1$1$1$2
X$28 VDD vias_gen$15$2$1$1$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$1$1$1$2

.SUBCKT rovcel2_LVT$1$1$1$1$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$1$1$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$1$1$1$2
X$3 IN GND OUT nfet$4$1$1$1$1$1$2
X$4 GND vias_gen$17$1$1$1$1$1$1$2
X$5 GND vias_gen$15$1$1$1$1$1$1$2
X$6 GND vias_gen$17$1$1$1$1$1$1$2
X$7 IN OUT GND nfet$4$1$1$1$1$1$2
X$8 OUT vias_gen$12$1$1$1$1$1$1$2
X$9 OUT vias_gen$8$1$1$1$1$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$1$1$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$1$1$1$2
X$12 OUT vias_gen$8$1$1$1$1$1$1$2
X$13 OUT vias_gen$12$1$1$1$1$1$1$2
X$14 OUT vias_gen$16$1$1$1$1$1$1$2
X$15 OUT vias_gen$16$1$1$1$1$1$1$2
X$16 IN OUT VDD VDD pfet$4$1$1$1$1$1$1$2
X$17 OUT vias_gen$13$1$1$1$1$1$1$2
X$18 IN VDD OUT VDD pfet$4$1$1$1$1$1$1$2
X$19 OUT vias_gen$13$1$1$1$1$1$1$2
X$20 IN VDD OUT VDD pfet$4$1$1$1$1$1$1$2
X$21 IN OUT VDD VDD pfet$4$1$1$1$1$1$1$2
X$22 IN vias_gen$14$1$1$1$1$1$1$2
X$23 IN vias_gen$14$1$1$1$1$1$1$2
X$24 IN vias_gen$14$1$1$1$1$1$1$2
X$25 IN vias_gen$14$1$1$1$1$1$1$2
X$26 VDD vias_gen$17$1$1$1$1$1$1$2
X$27 VDD vias_gen$15$1$1$1$1$1$1$2
X$28 VDD vias_gen$17$1$1$1$1$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$1$1$1$2

.SUBCKT rovcel2_LVT$3$1$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$1$1$1$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$1$1$1$2
X$3 IN OUT GND nfet$6$1$1$1$2
X$4 IN GND OUT nfet$6$1$1$1$2
X$5 GND vias_gen$17$3$1$1$1$2
X$6 GND vias_gen$17$3$1$1$1$2
X$7 GND vias_gen$15$3$1$1$1$2
X$8 OUT vias_gen$12$3$1$1$1$2
X$9 OUT vias_gen$8$3$1$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$3$1$1$1$2
X$11 VDD VDD \$28 OUT pfet$5$3$1$1$1$2
X$12 OUT vias_gen$8$3$1$1$1$2
X$13 OUT vias_gen$12$3$1$1$1$2
X$14 IN OUT VDD VDD pfet$4$3$1$1$1$2
X$15 IN VDD OUT VDD pfet$4$3$1$1$1$2
X$16 OUT vias_gen$13$3$1$1$1$2
X$17 IN VDD OUT VDD pfet$4$3$1$1$1$2
X$18 OUT vias_gen$13$3$1$1$1$2
X$19 IN OUT VDD VDD pfet$4$3$1$1$1$2
X$20 OUT vias_gen$16$3$1$1$1$2
X$21 OUT vias_gen$16$3$1$1$1$2
X$22 IN vias_gen$14$3$1$1$1$2
X$23 IN vias_gen$14$3$1$1$1$2
X$24 IN vias_gen$14$3$1$1$1$2
X$25 IN vias_gen$14$3$1$1$1$2
X$26 VDD vias_gen$17$3$1$1$1$2
X$27 VDD vias_gen$17$3$1$1$1$2
X$28 VDD vias_gen$15$3$1$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$1$1$1$2

.SUBCKT rovcel2_LVT$1$2$1$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$1$1$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$1$1$1$2
X$3 IN GND OUT nfet$4$2$1$1$1$2
X$4 GND vias_gen$17$1$2$1$1$1$2
X$5 GND vias_gen$15$1$2$1$1$1$2
X$6 GND vias_gen$17$1$2$1$1$1$2
X$7 IN OUT GND nfet$4$2$1$1$1$2
X$8 OUT vias_gen$12$1$2$1$1$1$2
X$9 OUT vias_gen$8$1$2$1$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$2$1$1$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$2$1$1$1$2
X$12 OUT vias_gen$8$1$2$1$1$1$2
X$13 OUT vias_gen$12$1$2$1$1$1$2
X$14 OUT vias_gen$16$1$2$1$1$1$2
X$15 OUT vias_gen$16$1$2$1$1$1$2
X$16 IN OUT VDD VDD pfet$4$1$2$1$1$1$2
X$17 OUT vias_gen$13$1$2$1$1$1$2
X$18 IN VDD OUT VDD pfet$4$1$2$1$1$1$2
X$19 OUT vias_gen$13$1$2$1$1$1$2
X$20 IN VDD OUT VDD pfet$4$1$2$1$1$1$2
X$21 IN OUT VDD VDD pfet$4$1$2$1$1$1$2
X$22 IN vias_gen$14$1$2$1$1$1$2
X$23 IN vias_gen$14$1$2$1$1$1$2
X$24 IN vias_gen$14$1$2$1$1$1$2
X$25 IN vias_gen$14$1$2$1$1$1$2
X$26 VDD vias_gen$17$1$2$1$1$1$2
X$27 VDD vias_gen$15$1$2$1$1$1$2
X$28 VDD vias_gen$17$1$2$1$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$1$1$1$2

.SUBCKT rovcel2_LVT$2$2$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$2$1$1$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$2$1$1$2
X$3 IN OUT GND nfet$5$2$1$1$2
X$4 IN GND OUT nfet$5$2$1$1$2
X$5 GND vias_gen$17$2$2$1$1$2
X$6 GND vias_gen$17$2$2$1$1$2
X$7 GND vias_gen$15$2$2$1$1$2
X$8 OUT vias_gen$12$2$2$1$1$2
X$9 OUT vias_gen$8$2$2$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$2$2$1$1$2
X$11 VDD VDD \$28 OUT pfet$5$2$2$1$1$2
X$12 OUT vias_gen$8$2$2$1$1$2
X$13 OUT vias_gen$12$2$2$1$1$2
X$14 IN OUT VDD VDD pfet$4$2$2$1$1$2
X$15 IN VDD OUT VDD pfet$4$2$2$1$1$2
X$16 OUT vias_gen$13$2$2$1$1$2
X$17 IN VDD OUT VDD pfet$4$2$2$1$1$2
X$18 OUT vias_gen$13$2$2$1$1$2
X$19 IN OUT VDD VDD pfet$4$2$2$1$1$2
X$20 OUT vias_gen$16$2$2$1$1$2
X$21 OUT vias_gen$16$2$2$1$1$2
X$22 IN vias_gen$14$2$2$1$1$2
X$23 IN vias_gen$14$2$2$1$1$2
X$24 IN vias_gen$14$2$2$1$1$2
X$25 IN vias_gen$14$2$2$1$1$2
X$26 VDD vias_gen$17$2$2$1$1$2
X$27 VDD vias_gen$17$2$2$1$1$2
X$28 VDD vias_gen$15$2$2$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$2$1$1$2

.SUBCKT rovcel2_LVT$1$1$2$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$2$1$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$2$1$1$2
X$3 IN GND OUT nfet$4$1$2$1$1$2
X$4 GND vias_gen$17$1$1$2$1$1$2
X$5 GND vias_gen$15$1$1$2$1$1$2
X$6 GND vias_gen$17$1$1$2$1$1$2
X$7 IN OUT GND nfet$4$1$2$1$1$2
X$8 OUT vias_gen$12$1$1$2$1$1$2
X$9 OUT vias_gen$8$1$1$2$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$1$2$1$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$1$2$1$1$2
X$12 OUT vias_gen$8$1$1$2$1$1$2
X$13 OUT vias_gen$12$1$1$2$1$1$2
X$14 OUT vias_gen$16$1$1$2$1$1$2
X$15 OUT vias_gen$16$1$1$2$1$1$2
X$16 IN OUT VDD VDD pfet$4$1$1$2$1$1$2
X$17 OUT vias_gen$13$1$1$2$1$1$2
X$18 IN VDD OUT VDD pfet$4$1$1$2$1$1$2
X$19 OUT vias_gen$13$1$1$2$1$1$2
X$20 IN VDD OUT VDD pfet$4$1$1$2$1$1$2
X$21 IN OUT VDD VDD pfet$4$1$1$2$1$1$2
X$22 IN vias_gen$14$1$1$2$1$1$2
X$23 IN vias_gen$14$1$1$2$1$1$2
X$24 IN vias_gen$14$1$1$2$1$1$2
X$25 IN vias_gen$14$1$1$2$1$1$2
X$26 VDD vias_gen$17$1$1$2$1$1$2
X$27 VDD vias_gen$15$1$1$2$1$1$2
X$28 VDD vias_gen$17$1$1$2$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$2$1$1$2

.SUBCKT rovcel2_LVT$2$1$2$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$2$1$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$2$1$2
X$3 IN OUT GND nfet$5$1$2$1$2
X$4 IN GND OUT nfet$5$1$2$1$2
X$5 GND vias_gen$17$2$1$2$1$2
X$6 GND vias_gen$17$2$1$2$1$2
X$7 GND vias_gen$15$2$1$2$1$2
X$8 OUT vias_gen$12$2$1$2$1$2
X$9 OUT vias_gen$8$2$1$2$1$2
X$10 VDD VDD \$25 OUT pfet$5$2$1$2$1$2
X$11 VDD VDD \$28 OUT pfet$5$2$1$2$1$2
X$12 OUT vias_gen$8$2$1$2$1$2
X$13 OUT vias_gen$12$2$1$2$1$2
X$14 IN OUT VDD VDD pfet$4$2$1$2$1$2
X$15 IN VDD OUT VDD pfet$4$2$1$2$1$2
X$16 OUT vias_gen$13$2$1$2$1$2
X$17 IN VDD OUT VDD pfet$4$2$1$2$1$2
X$18 OUT vias_gen$13$2$1$2$1$2
X$19 IN OUT VDD VDD pfet$4$2$1$2$1$2
X$20 OUT vias_gen$16$2$1$2$1$2
X$21 OUT vias_gen$16$2$1$2$1$2
X$22 IN vias_gen$14$2$1$2$1$2
X$23 IN vias_gen$14$2$1$2$1$2
X$24 IN vias_gen$14$2$1$2$1$2
X$25 IN vias_gen$14$2$1$2$1$2
X$26 VDD vias_gen$17$2$1$2$1$2
X$27 VDD vias_gen$17$2$1$2$1$2
X$28 VDD vias_gen$15$2$1$2$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$2$1$2

.SUBCKT rovcel2_LVT$1$1$1$2$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$2$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$2$1$2
X$3 IN GND OUT nfet$4$1$1$2$1$2
X$4 GND vias_gen$17$1$1$1$2$1$2
X$5 GND vias_gen$15$1$1$1$2$1$2
X$6 GND vias_gen$17$1$1$1$2$1$2
X$7 IN OUT GND nfet$4$1$1$2$1$2
X$8 OUT vias_gen$12$1$1$1$2$1$2
X$9 OUT vias_gen$8$1$1$1$2$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$2$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$2$1$2
X$12 OUT vias_gen$8$1$1$1$2$1$2
X$13 OUT vias_gen$12$1$1$1$2$1$2
X$14 OUT vias_gen$16$1$1$1$2$1$2
X$15 OUT vias_gen$16$1$1$1$2$1$2
X$16 IN OUT VDD VDD pfet$4$1$1$1$2$1$2
X$17 OUT vias_gen$13$1$1$1$2$1$2
X$18 IN VDD OUT VDD pfet$4$1$1$1$2$1$2
X$19 OUT vias_gen$13$1$1$1$2$1$2
X$20 IN VDD OUT VDD pfet$4$1$1$1$2$1$2
X$21 IN OUT VDD VDD pfet$4$1$1$1$2$1$2
X$22 IN vias_gen$14$1$1$1$2$1$2
X$23 IN vias_gen$14$1$1$1$2$1$2
X$24 IN vias_gen$14$1$1$1$2$1$2
X$25 IN vias_gen$14$1$1$1$2$1$2
X$26 VDD vias_gen$17$1$1$1$2$1$2
X$27 VDD vias_gen$15$1$1$1$2$1$2
X$28 VDD vias_gen$17$1$1$1$2$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$2$1$2

.SUBCKT rovcel2_LVT$3$2$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$2$1$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$2$1$2
X$3 IN OUT GND nfet$6$2$1$2
X$4 IN GND OUT nfet$6$2$1$2
X$5 GND vias_gen$17$3$2$1$2
X$6 GND vias_gen$17$3$2$1$2
X$7 GND vias_gen$15$3$2$1$2
X$8 OUT vias_gen$12$3$2$1$2
X$9 OUT vias_gen$8$3$2$1$2
X$10 VDD VDD \$25 OUT pfet$5$3$2$1$2
X$11 VDD VDD \$28 OUT pfet$5$3$2$1$2
X$12 OUT vias_gen$8$3$2$1$2
X$13 OUT vias_gen$12$3$2$1$2
X$14 IN OUT VDD VDD pfet$4$3$2$1$2
X$15 IN VDD OUT VDD pfet$4$3$2$1$2
X$16 OUT vias_gen$13$3$2$1$2
X$17 IN VDD OUT VDD pfet$4$3$2$1$2
X$18 OUT vias_gen$13$3$2$1$2
X$19 IN OUT VDD VDD pfet$4$3$2$1$2
X$20 OUT vias_gen$16$3$2$1$2
X$21 OUT vias_gen$16$3$2$1$2
X$22 IN vias_gen$14$3$2$1$2
X$23 IN vias_gen$14$3$2$1$2
X$24 IN vias_gen$14$3$2$1$2
X$25 IN vias_gen$14$3$2$1$2
X$26 VDD vias_gen$17$3$2$1$2
X$27 VDD vias_gen$17$3$2$1$2
X$28 VDD vias_gen$15$3$2$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$2$1$2

.SUBCKT rovcel2_LVT$1$2$2$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$2$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$2$1$2
X$3 IN GND OUT nfet$4$2$2$1$2
X$4 GND vias_gen$17$1$2$2$1$2
X$5 GND vias_gen$15$1$2$2$1$2
X$6 GND vias_gen$17$1$2$2$1$2
X$7 IN OUT GND nfet$4$2$2$1$2
X$8 OUT vias_gen$12$1$2$2$1$2
X$9 OUT vias_gen$8$1$2$2$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$2$2$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$2$2$1$2
X$12 OUT vias_gen$8$1$2$2$1$2
X$13 OUT vias_gen$12$1$2$2$1$2
X$14 OUT vias_gen$16$1$2$2$1$2
X$15 OUT vias_gen$16$1$2$2$1$2
X$16 IN OUT VDD VDD pfet$4$1$2$2$1$2
X$17 OUT vias_gen$13$1$2$2$1$2
X$18 IN VDD OUT VDD pfet$4$1$2$2$1$2
X$19 OUT vias_gen$13$1$2$2$1$2
X$20 IN VDD OUT VDD pfet$4$1$2$2$1$2
X$21 IN OUT VDD VDD pfet$4$1$2$2$1$2
X$22 IN vias_gen$14$1$2$2$1$2
X$23 IN vias_gen$14$1$2$2$1$2
X$24 IN vias_gen$14$1$2$2$1$2
X$25 IN vias_gen$14$1$2$2$1$2
X$26 VDD vias_gen$17$1$2$2$1$2
X$27 VDD vias_gen$15$1$2$2$1$2
X$28 VDD vias_gen$17$1$2$2$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$2$1$2

.SUBCKT rovcel2_LVT$2$1$1$1$3 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$1$1$3
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$1$1$3
X$3 IN OUT GND nfet$5$1$1$1$3
X$4 IN GND OUT nfet$5$1$1$1$3
X$5 GND vias_gen$17$2$1$1$1$3
X$6 GND vias_gen$17$2$1$1$1$3
X$7 GND vias_gen$15$2$1$1$1$3
X$8 OUT vias_gen$12$2$1$1$1$3
X$9 OUT vias_gen$8$2$1$1$1$3
X$10 VDD VDD \$25 OUT pfet$5$2$1$1$1$3
X$11 VDD VDD \$28 OUT pfet$5$2$1$1$1$3
X$12 OUT vias_gen$8$2$1$1$1$3
X$13 OUT vias_gen$12$2$1$1$1$3
X$14 IN OUT VDD VDD pfet$4$2$1$1$1$3
X$15 IN VDD OUT VDD pfet$4$2$1$1$1$3
X$16 OUT vias_gen$13$2$1$1$1$3
X$17 IN VDD OUT VDD pfet$4$2$1$1$1$3
X$18 OUT vias_gen$13$2$1$1$1$3
X$19 IN OUT VDD VDD pfet$4$2$1$1$1$3
X$20 OUT vias_gen$16$2$1$1$1$3
X$21 OUT vias_gen$16$2$1$1$1$3
X$22 IN vias_gen$14$2$1$1$1$3
X$23 IN vias_gen$14$2$1$1$1$3
X$24 IN vias_gen$14$2$1$1$1$3
X$25 IN vias_gen$14$2$1$1$1$3
X$26 VDD vias_gen$17$2$1$1$1$3
X$27 VDD vias_gen$17$2$1$1$1$3
X$28 VDD vias_gen$15$2$1$1$1$3
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$1$1$3

.SUBCKT rovcel2_LVT$1$1$1$1$1$3 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$1$1$3
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$1$1$3
X$3 IN GND OUT nfet$4$1$1$1$1$3
X$4 GND vias_gen$17$1$1$1$1$1$3
X$5 GND vias_gen$15$1$1$1$1$1$3
X$6 GND vias_gen$17$1$1$1$1$1$3
X$7 IN OUT GND nfet$4$1$1$1$1$3
X$8 OUT vias_gen$12$1$1$1$1$1$3
X$9 OUT vias_gen$8$1$1$1$1$1$3
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$1$1$3
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$1$1$3
X$12 OUT vias_gen$8$1$1$1$1$1$3
X$13 OUT vias_gen$12$1$1$1$1$1$3
X$14 OUT vias_gen$16$1$1$1$1$1$3
X$15 OUT vias_gen$16$1$1$1$1$1$3
X$16 IN OUT VDD VDD pfet$4$1$1$1$1$1$3
X$17 OUT vias_gen$13$1$1$1$1$1$3
X$18 IN VDD OUT VDD pfet$4$1$1$1$1$1$3
X$19 OUT vias_gen$13$1$1$1$1$1$3
X$20 IN VDD OUT VDD pfet$4$1$1$1$1$1$3
X$21 IN OUT VDD VDD pfet$4$1$1$1$1$1$3
X$22 IN vias_gen$14$1$1$1$1$1$3
X$23 IN vias_gen$14$1$1$1$1$1$3
X$24 IN vias_gen$14$1$1$1$1$1$3
X$25 IN vias_gen$14$1$1$1$1$1$3
X$26 VDD vias_gen$17$1$1$1$1$1$3
X$27 VDD vias_gen$15$1$1$1$1$1$3
X$28 VDD vias_gen$17$1$1$1$1$1$3
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$1$1$3

.SUBCKT rovcel2_LVT$3$1$1$3 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$1$1$3
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$1$1$3
X$3 IN OUT GND nfet$6$1$1$3
X$4 IN GND OUT nfet$6$1$1$3
X$5 GND vias_gen$17$3$1$1$3
X$6 GND vias_gen$17$3$1$1$3
X$7 GND vias_gen$15$3$1$1$3
X$8 OUT vias_gen$12$3$1$1$3
X$9 OUT vias_gen$8$3$1$1$3
X$10 VDD VDD \$25 OUT pfet$5$3$1$1$3
X$11 VDD VDD \$28 OUT pfet$5$3$1$1$3
X$12 OUT vias_gen$8$3$1$1$3
X$13 OUT vias_gen$12$3$1$1$3
X$14 IN OUT VDD VDD pfet$4$3$1$1$3
X$15 IN VDD OUT VDD pfet$4$3$1$1$3
X$16 OUT vias_gen$13$3$1$1$3
X$17 IN VDD OUT VDD pfet$4$3$1$1$3
X$18 OUT vias_gen$13$3$1$1$3
X$19 IN OUT VDD VDD pfet$4$3$1$1$3
X$20 OUT vias_gen$16$3$1$1$3
X$21 OUT vias_gen$16$3$1$1$3
X$22 IN vias_gen$14$3$1$1$3
X$23 IN vias_gen$14$3$1$1$3
X$24 IN vias_gen$14$3$1$1$3
X$25 IN vias_gen$14$3$1$1$3
X$26 VDD vias_gen$17$3$1$1$3
X$27 VDD vias_gen$17$3$1$1$3
X$28 VDD vias_gen$15$3$1$1$3
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$1$1$3

.SUBCKT rovcel2_LVT$1$2$1$1$3 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$1$1$3
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$1$1$3
X$3 IN GND OUT nfet$4$2$1$1$3
X$4 GND vias_gen$17$1$2$1$1$3
X$5 GND vias_gen$15$1$2$1$1$3
X$6 GND vias_gen$17$1$2$1$1$3
X$7 IN OUT GND nfet$4$2$1$1$3
X$8 OUT vias_gen$12$1$2$1$1$3
X$9 OUT vias_gen$8$1$2$1$1$3
X$10 VDD VDD \$25 OUT pfet$5$1$2$1$1$3
X$11 VDD VDD \$27 OUT pfet$5$1$2$1$1$3
X$12 OUT vias_gen$8$1$2$1$1$3
X$13 OUT vias_gen$12$1$2$1$1$3
X$14 OUT vias_gen$16$1$2$1$1$3
X$15 OUT vias_gen$16$1$2$1$1$3
X$16 IN OUT VDD VDD pfet$4$1$2$1$1$3
X$17 OUT vias_gen$13$1$2$1$1$3
X$18 IN VDD OUT VDD pfet$4$1$2$1$1$3
X$19 OUT vias_gen$13$1$2$1$1$3
X$20 IN VDD OUT VDD pfet$4$1$2$1$1$3
X$21 IN OUT VDD VDD pfet$4$1$2$1$1$3
X$22 IN vias_gen$14$1$2$1$1$3
X$23 IN vias_gen$14$1$2$1$1$3
X$24 IN vias_gen$14$1$2$1$1$3
X$25 IN vias_gen$14$1$2$1$1$3
X$26 VDD vias_gen$17$1$2$1$1$3
X$27 VDD vias_gen$15$1$2$1$1$3
X$28 VDD vias_gen$17$1$2$1$1$3
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$1$1$3

.SUBCKT rovcel2_LVT$2$1$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$1$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$1$1$1$1
X$3 IN OUT GND nfet$5$1$1$1$1$1
X$4 IN GND OUT nfet$5$1$1$1$1$1
X$5 GND vias_gen$17$2$1$1$1$1$1
X$6 GND vias_gen$17$2$1$1$1$1$1
X$7 GND vias_gen$15$2$1$1$1$1$1
X$8 OUT vias_gen$12$2$1$1$1$1$1
X$9 OUT vias_gen$8$2$1$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$2$1$1$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$2$1$1$1$1$1
X$12 OUT vias_gen$8$2$1$1$1$1$1
X$13 OUT vias_gen$12$2$1$1$1$1$1
X$14 IN OUT VDD VDD pfet$4$2$1$1$1$1$1
X$15 IN VDD OUT VDD pfet$4$2$1$1$1$1$1
X$16 OUT vias_gen$13$2$1$1$1$1$1
X$17 IN VDD OUT VDD pfet$4$2$1$1$1$1$1
X$18 OUT vias_gen$13$2$1$1$1$1$1
X$19 IN OUT VDD VDD pfet$4$2$1$1$1$1$1
X$20 OUT vias_gen$16$2$1$1$1$1$1
X$21 OUT vias_gen$16$2$1$1$1$1$1
X$22 IN vias_gen$14$2$1$1$1$1$1
X$23 IN vias_gen$14$2$1$1$1$1$1
X$24 IN vias_gen$14$2$1$1$1$1$1
X$25 IN vias_gen$14$2$1$1$1$1$1
X$26 VDD vias_gen$17$2$1$1$1$1$1
X$27 VDD vias_gen$17$2$1$1$1$1$1
X$28 VDD vias_gen$15$2$1$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$1$1$1$1

.SUBCKT rovcel2_LVT$1$1$1$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$1$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$1$1$1$1
X$3 IN GND OUT nfet$4$1$1$1$1$1$1
X$4 GND vias_gen$17$1$1$1$1$1$1$1
X$5 GND vias_gen$15$1$1$1$1$1$1$1
X$6 GND vias_gen$17$1$1$1$1$1$1$1
X$7 IN OUT GND nfet$4$1$1$1$1$1$1
X$8 OUT vias_gen$12$1$1$1$1$1$1$1
X$9 OUT vias_gen$8$1$1$1$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$1$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$1$1$1$1
X$12 OUT vias_gen$8$1$1$1$1$1$1$1
X$13 OUT vias_gen$12$1$1$1$1$1$1$1
X$14 OUT vias_gen$16$1$1$1$1$1$1$1
X$15 OUT vias_gen$16$1$1$1$1$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$1$1$1$1$1
X$17 OUT vias_gen$13$1$1$1$1$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$1$1$1$1$1
X$19 OUT vias_gen$13$1$1$1$1$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$1$1$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$1$1$1$1$1
X$22 IN vias_gen$14$1$1$1$1$1$1$1
X$23 IN vias_gen$14$1$1$1$1$1$1$1
X$24 IN vias_gen$14$1$1$1$1$1$1$1
X$25 IN vias_gen$14$1$1$1$1$1$1$1
X$26 VDD vias_gen$17$1$1$1$1$1$1$1
X$27 VDD vias_gen$15$1$1$1$1$1$1$1
X$28 VDD vias_gen$17$1$1$1$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$1$1$1$1

.SUBCKT rovcel2_LVT$3$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$1$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$1$1$1$1
X$3 IN OUT GND nfet$6$1$1$1$1
X$4 IN GND OUT nfet$6$1$1$1$1
X$5 GND vias_gen$17$3$1$1$1$1
X$6 GND vias_gen$17$3$1$1$1$1
X$7 GND vias_gen$15$3$1$1$1$1
X$8 OUT vias_gen$12$3$1$1$1$1
X$9 OUT vias_gen$8$3$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$3$1$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$3$1$1$1$1
X$12 OUT vias_gen$8$3$1$1$1$1
X$13 OUT vias_gen$12$3$1$1$1$1
X$14 IN OUT VDD VDD pfet$4$3$1$1$1$1
X$15 IN VDD OUT VDD pfet$4$3$1$1$1$1
X$16 OUT vias_gen$13$3$1$1$1$1
X$17 IN VDD OUT VDD pfet$4$3$1$1$1$1
X$18 OUT vias_gen$13$3$1$1$1$1
X$19 IN OUT VDD VDD pfet$4$3$1$1$1$1
X$20 OUT vias_gen$16$3$1$1$1$1
X$21 OUT vias_gen$16$3$1$1$1$1
X$22 IN vias_gen$14$3$1$1$1$1
X$23 IN vias_gen$14$3$1$1$1$1
X$24 IN vias_gen$14$3$1$1$1$1
X$25 IN vias_gen$14$3$1$1$1$1
X$26 VDD vias_gen$17$3$1$1$1$1
X$27 VDD vias_gen$17$3$1$1$1$1
X$28 VDD vias_gen$15$3$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$1$1$1$1

.SUBCKT rovcel2_LVT$1$2$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$1$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$1$1$1$1
X$3 IN GND OUT nfet$4$2$1$1$1$1
X$4 GND vias_gen$17$1$2$1$1$1$1
X$5 GND vias_gen$15$1$2$1$1$1$1
X$6 GND vias_gen$17$1$2$1$1$1$1
X$7 IN OUT GND nfet$4$2$1$1$1$1
X$8 OUT vias_gen$12$1$2$1$1$1$1
X$9 OUT vias_gen$8$1$2$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$2$1$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$2$1$1$1$1
X$12 OUT vias_gen$8$1$2$1$1$1$1
X$13 OUT vias_gen$12$1$2$1$1$1$1
X$14 OUT vias_gen$16$1$2$1$1$1$1
X$15 OUT vias_gen$16$1$2$1$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$2$1$1$1$1
X$17 OUT vias_gen$13$1$2$1$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$2$1$1$1$1
X$19 OUT vias_gen$13$1$2$1$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$2$1$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$2$1$1$1$1
X$22 IN vias_gen$14$1$2$1$1$1$1
X$23 IN vias_gen$14$1$2$1$1$1$1
X$24 IN vias_gen$14$1$2$1$1$1$1
X$25 IN vias_gen$14$1$2$1$1$1$1
X$26 VDD vias_gen$17$1$2$1$1$1$1
X$27 VDD vias_gen$15$1$2$1$1$1$1
X$28 VDD vias_gen$17$1$2$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$1$1$1$1

.SUBCKT rovcel2_LVT$2$2$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$2$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$2$1$1$1
X$3 IN OUT GND nfet$5$2$1$1$1
X$4 IN GND OUT nfet$5$2$1$1$1
X$5 GND vias_gen$17$2$2$1$1$1
X$6 GND vias_gen$17$2$2$1$1$1
X$7 GND vias_gen$15$2$2$1$1$1
X$8 OUT vias_gen$12$2$2$1$1$1
X$9 OUT vias_gen$8$2$2$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$2$2$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$2$2$1$1$1
X$12 OUT vias_gen$8$2$2$1$1$1
X$13 OUT vias_gen$12$2$2$1$1$1
X$14 IN OUT VDD VDD pfet$4$2$2$1$1$1
X$15 IN VDD OUT VDD pfet$4$2$2$1$1$1
X$16 OUT vias_gen$13$2$2$1$1$1
X$17 IN VDD OUT VDD pfet$4$2$2$1$1$1
X$18 OUT vias_gen$13$2$2$1$1$1
X$19 IN OUT VDD VDD pfet$4$2$2$1$1$1
X$20 OUT vias_gen$16$2$2$1$1$1
X$21 OUT vias_gen$16$2$2$1$1$1
X$22 IN vias_gen$14$2$2$1$1$1
X$23 IN vias_gen$14$2$2$1$1$1
X$24 IN vias_gen$14$2$2$1$1$1
X$25 IN vias_gen$14$2$2$1$1$1
X$26 VDD vias_gen$17$2$2$1$1$1
X$27 VDD vias_gen$17$2$2$1$1$1
X$28 VDD vias_gen$15$2$2$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$2$1$1$1

.SUBCKT rovcel2_LVT$1$1$2$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$2$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$2$1$1$1
X$3 IN GND OUT nfet$4$1$2$1$1$1
X$4 GND vias_gen$17$1$1$2$1$1$1
X$5 GND vias_gen$15$1$1$2$1$1$1
X$6 GND vias_gen$17$1$1$2$1$1$1
X$7 IN OUT GND nfet$4$1$2$1$1$1
X$8 OUT vias_gen$12$1$1$2$1$1$1
X$9 OUT vias_gen$8$1$1$2$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$2$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$2$1$1$1
X$12 OUT vias_gen$8$1$1$2$1$1$1
X$13 OUT vias_gen$12$1$1$2$1$1$1
X$14 OUT vias_gen$16$1$1$2$1$1$1
X$15 OUT vias_gen$16$1$1$2$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$2$1$1$1
X$17 OUT vias_gen$13$1$1$2$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$2$1$1$1
X$19 OUT vias_gen$13$1$1$2$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$2$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$2$1$1$1
X$22 IN vias_gen$14$1$1$2$1$1$1
X$23 IN vias_gen$14$1$1$2$1$1$1
X$24 IN vias_gen$14$1$1$2$1$1$1
X$25 IN vias_gen$14$1$1$2$1$1$1
X$26 VDD vias_gen$17$1$1$2$1$1$1
X$27 VDD vias_gen$15$1$1$2$1$1$1
X$28 VDD vias_gen$17$1$1$2$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$2$1$1$1

.SUBCKT rovcel2_LVT$2$1$2$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$2$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$2$1$1
X$3 IN OUT GND nfet$5$1$2$1$1
X$4 IN GND OUT nfet$5$1$2$1$1
X$5 GND vias_gen$17$2$1$2$1$1
X$6 GND vias_gen$17$2$1$2$1$1
X$7 GND vias_gen$15$2$1$2$1$1
X$8 OUT vias_gen$12$2$1$2$1$1
X$9 OUT vias_gen$8$2$1$2$1$1
X$10 VDD VDD \$25 OUT pfet$5$2$1$2$1$1
X$11 VDD VDD \$28 OUT pfet$5$2$1$2$1$1
X$12 OUT vias_gen$8$2$1$2$1$1
X$13 OUT vias_gen$12$2$1$2$1$1
X$14 IN OUT VDD VDD pfet$4$2$1$2$1$1
X$15 IN VDD OUT VDD pfet$4$2$1$2$1$1
X$16 OUT vias_gen$13$2$1$2$1$1
X$17 IN VDD OUT VDD pfet$4$2$1$2$1$1
X$18 OUT vias_gen$13$2$1$2$1$1
X$19 IN OUT VDD VDD pfet$4$2$1$2$1$1
X$20 OUT vias_gen$16$2$1$2$1$1
X$21 OUT vias_gen$16$2$1$2$1$1
X$22 IN vias_gen$14$2$1$2$1$1
X$23 IN vias_gen$14$2$1$2$1$1
X$24 IN vias_gen$14$2$1$2$1$1
X$25 IN vias_gen$14$2$1$2$1$1
X$26 VDD vias_gen$17$2$1$2$1$1
X$27 VDD vias_gen$17$2$1$2$1$1
X$28 VDD vias_gen$15$2$1$2$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$2$1$1

.SUBCKT rovcel2_LVT$1$1$1$2$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$2$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$2$1$1
X$3 IN GND OUT nfet$4$1$1$2$1$1
X$4 GND vias_gen$17$1$1$1$2$1$1
X$5 GND vias_gen$15$1$1$1$2$1$1
X$6 GND vias_gen$17$1$1$1$2$1$1
X$7 IN OUT GND nfet$4$1$1$2$1$1
X$8 OUT vias_gen$12$1$1$1$2$1$1
X$9 OUT vias_gen$8$1$1$1$2$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$2$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$2$1$1
X$12 OUT vias_gen$8$1$1$1$2$1$1
X$13 OUT vias_gen$12$1$1$1$2$1$1
X$14 OUT vias_gen$16$1$1$1$2$1$1
X$15 OUT vias_gen$16$1$1$1$2$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$1$2$1$1
X$17 OUT vias_gen$13$1$1$1$2$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$1$2$1$1
X$19 OUT vias_gen$13$1$1$1$2$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$1$2$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$1$2$1$1
X$22 IN vias_gen$14$1$1$1$2$1$1
X$23 IN vias_gen$14$1$1$1$2$1$1
X$24 IN vias_gen$14$1$1$1$2$1$1
X$25 IN vias_gen$14$1$1$1$2$1$1
X$26 VDD vias_gen$17$1$1$1$2$1$1
X$27 VDD vias_gen$15$1$1$1$2$1$1
X$28 VDD vias_gen$17$1$1$1$2$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$2$1$1

.SUBCKT rovcel2_LVT$3$2$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$2$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$2$1$1
X$3 IN OUT GND nfet$6$2$1$1
X$4 IN GND OUT nfet$6$2$1$1
X$5 GND vias_gen$17$3$2$1$1
X$6 GND vias_gen$17$3$2$1$1
X$7 GND vias_gen$15$3$2$1$1
X$8 OUT vias_gen$12$3$2$1$1
X$9 OUT vias_gen$8$3$2$1$1
X$10 VDD VDD \$25 OUT pfet$5$3$2$1$1
X$11 VDD VDD \$28 OUT pfet$5$3$2$1$1
X$12 OUT vias_gen$8$3$2$1$1
X$13 OUT vias_gen$12$3$2$1$1
X$14 IN OUT VDD VDD pfet$4$3$2$1$1
X$15 IN VDD OUT VDD pfet$4$3$2$1$1
X$16 OUT vias_gen$13$3$2$1$1
X$17 IN VDD OUT VDD pfet$4$3$2$1$1
X$18 OUT vias_gen$13$3$2$1$1
X$19 IN OUT VDD VDD pfet$4$3$2$1$1
X$20 OUT vias_gen$16$3$2$1$1
X$21 OUT vias_gen$16$3$2$1$1
X$22 IN vias_gen$14$3$2$1$1
X$23 IN vias_gen$14$3$2$1$1
X$24 IN vias_gen$14$3$2$1$1
X$25 IN vias_gen$14$3$2$1$1
X$26 VDD vias_gen$17$3$2$1$1
X$27 VDD vias_gen$17$3$2$1$1
X$28 VDD vias_gen$15$3$2$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$2$1$1

.SUBCKT rovcel2_LVT$1$2$2$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$2$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$2$1$1
X$3 IN GND OUT nfet$4$2$2$1$1
X$4 GND vias_gen$17$1$2$2$1$1
X$5 GND vias_gen$15$1$2$2$1$1
X$6 GND vias_gen$17$1$2$2$1$1
X$7 IN OUT GND nfet$4$2$2$1$1
X$8 OUT vias_gen$12$1$2$2$1$1
X$9 OUT vias_gen$8$1$2$2$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$2$2$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$2$2$1$1
X$12 OUT vias_gen$8$1$2$2$1$1
X$13 OUT vias_gen$12$1$2$2$1$1
X$14 OUT vias_gen$16$1$2$2$1$1
X$15 OUT vias_gen$16$1$2$2$1$1
X$16 IN OUT VDD VDD pfet$4$1$2$2$1$1
X$17 OUT vias_gen$13$1$2$2$1$1
X$18 IN VDD OUT VDD pfet$4$1$2$2$1$1
X$19 OUT vias_gen$13$1$2$2$1$1
X$20 IN VDD OUT VDD pfet$4$1$2$2$1$1
X$21 IN OUT VDD VDD pfet$4$1$2$2$1$1
X$22 IN vias_gen$14$1$2$2$1$1
X$23 IN vias_gen$14$1$2$2$1$1
X$24 IN vias_gen$14$1$2$2$1$1
X$25 IN vias_gen$14$1$2$2$1$1
X$26 VDD vias_gen$17$1$2$2$1$1
X$27 VDD vias_gen$15$1$2$2$1$1
X$28 VDD vias_gen$17$1$2$2$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$2$1$1

.SUBCKT rovcel2_LVT$2$1$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$1$1$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$1$1$2
X$3 IN OUT GND nfet$5$1$1$1$2
X$4 IN GND OUT nfet$5$1$1$1$2
X$5 GND vias_gen$17$2$1$1$1$2
X$6 GND vias_gen$17$2$1$1$1$2
X$7 GND vias_gen$15$2$1$1$1$2
X$8 OUT vias_gen$12$2$1$1$1$2
X$9 OUT vias_gen$8$2$1$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$2$1$1$1$2
X$11 VDD VDD \$28 OUT pfet$5$2$1$1$1$2
X$12 OUT vias_gen$8$2$1$1$1$2
X$13 OUT vias_gen$12$2$1$1$1$2
X$14 IN OUT VDD VDD pfet$4$2$1$1$1$2
X$15 IN VDD OUT VDD pfet$4$2$1$1$1$2
X$16 OUT vias_gen$13$2$1$1$1$2
X$17 IN VDD OUT VDD pfet$4$2$1$1$1$2
X$18 OUT vias_gen$13$2$1$1$1$2
X$19 IN OUT VDD VDD pfet$4$2$1$1$1$2
X$20 OUT vias_gen$16$2$1$1$1$2
X$21 OUT vias_gen$16$2$1$1$1$2
X$22 IN vias_gen$14$2$1$1$1$2
X$23 IN vias_gen$14$2$1$1$1$2
X$24 IN vias_gen$14$2$1$1$1$2
X$25 IN vias_gen$14$2$1$1$1$2
X$26 VDD vias_gen$17$2$1$1$1$2
X$27 VDD vias_gen$17$2$1$1$1$2
X$28 VDD vias_gen$15$2$1$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$1$1$2

.SUBCKT rovcel2_LVT$1$1$1$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$1$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$1$1$2
X$3 IN GND OUT nfet$4$1$1$1$1$2
X$4 GND vias_gen$17$1$1$1$1$1$2
X$5 GND vias_gen$15$1$1$1$1$1$2
X$6 GND vias_gen$17$1$1$1$1$1$2
X$7 IN OUT GND nfet$4$1$1$1$1$2
X$8 OUT vias_gen$12$1$1$1$1$1$2
X$9 OUT vias_gen$8$1$1$1$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$1$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$1$1$2
X$12 OUT vias_gen$8$1$1$1$1$1$2
X$13 OUT vias_gen$12$1$1$1$1$1$2
X$14 OUT vias_gen$16$1$1$1$1$1$2
X$15 OUT vias_gen$16$1$1$1$1$1$2
X$16 IN OUT VDD VDD pfet$4$1$1$1$1$1$2
X$17 OUT vias_gen$13$1$1$1$1$1$2
X$18 IN VDD OUT VDD pfet$4$1$1$1$1$1$2
X$19 OUT vias_gen$13$1$1$1$1$1$2
X$20 IN VDD OUT VDD pfet$4$1$1$1$1$1$2
X$21 IN OUT VDD VDD pfet$4$1$1$1$1$1$2
X$22 IN vias_gen$14$1$1$1$1$1$2
X$23 IN vias_gen$14$1$1$1$1$1$2
X$24 IN vias_gen$14$1$1$1$1$1$2
X$25 IN vias_gen$14$1$1$1$1$1$2
X$26 VDD vias_gen$17$1$1$1$1$1$2
X$27 VDD vias_gen$15$1$1$1$1$1$2
X$28 VDD vias_gen$17$1$1$1$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$1$1$2

.SUBCKT rovcel2_LVT$3$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$1$1$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$1$1$2
X$3 IN OUT GND nfet$6$1$1$2
X$4 IN GND OUT nfet$6$1$1$2
X$5 GND vias_gen$17$3$1$1$2
X$6 GND vias_gen$17$3$1$1$2
X$7 GND vias_gen$15$3$1$1$2
X$8 OUT vias_gen$12$3$1$1$2
X$9 OUT vias_gen$8$3$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$3$1$1$2
X$11 VDD VDD \$28 OUT pfet$5$3$1$1$2
X$12 OUT vias_gen$8$3$1$1$2
X$13 OUT vias_gen$12$3$1$1$2
X$14 IN OUT VDD VDD pfet$4$3$1$1$2
X$15 IN VDD OUT VDD pfet$4$3$1$1$2
X$16 OUT vias_gen$13$3$1$1$2
X$17 IN VDD OUT VDD pfet$4$3$1$1$2
X$18 OUT vias_gen$13$3$1$1$2
X$19 IN OUT VDD VDD pfet$4$3$1$1$2
X$20 OUT vias_gen$16$3$1$1$2
X$21 OUT vias_gen$16$3$1$1$2
X$22 IN vias_gen$14$3$1$1$2
X$23 IN vias_gen$14$3$1$1$2
X$24 IN vias_gen$14$3$1$1$2
X$25 IN vias_gen$14$3$1$1$2
X$26 VDD vias_gen$17$3$1$1$2
X$27 VDD vias_gen$17$3$1$1$2
X$28 VDD vias_gen$15$3$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$1$1$2

.SUBCKT rovcel2_LVT$1$2$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$1$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$1$1$2
X$3 IN GND OUT nfet$4$2$1$1$2
X$4 GND vias_gen$17$1$2$1$1$2
X$5 GND vias_gen$15$1$2$1$1$2
X$6 GND vias_gen$17$1$2$1$1$2
X$7 IN OUT GND nfet$4$2$1$1$2
X$8 OUT vias_gen$12$1$2$1$1$2
X$9 OUT vias_gen$8$1$2$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$2$1$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$2$1$1$2
X$12 OUT vias_gen$8$1$2$1$1$2
X$13 OUT vias_gen$12$1$2$1$1$2
X$14 OUT vias_gen$16$1$2$1$1$2
X$15 OUT vias_gen$16$1$2$1$1$2
X$16 IN OUT VDD VDD pfet$4$1$2$1$1$2
X$17 OUT vias_gen$13$1$2$1$1$2
X$18 IN VDD OUT VDD pfet$4$1$2$1$1$2
X$19 OUT vias_gen$13$1$2$1$1$2
X$20 IN VDD OUT VDD pfet$4$1$2$1$1$2
X$21 IN OUT VDD VDD pfet$4$1$2$1$1$2
X$22 IN vias_gen$14$1$2$1$1$2
X$23 IN vias_gen$14$1$2$1$1$2
X$24 IN vias_gen$14$1$2$1$1$2
X$25 IN vias_gen$14$1$2$1$1$2
X$26 VDD vias_gen$17$1$2$1$1$2
X$27 VDD vias_gen$15$1$2$1$1$2
X$28 VDD vias_gen$17$1$2$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$1$1$2

.SUBCKT rovcel2_LVT$2$2$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$2$1$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$2$1$2
X$3 IN OUT GND nfet$5$2$1$2
X$4 IN GND OUT nfet$5$2$1$2
X$5 GND vias_gen$17$2$2$1$2
X$6 GND vias_gen$17$2$2$1$2
X$7 GND vias_gen$15$2$2$1$2
X$8 OUT vias_gen$12$2$2$1$2
X$9 OUT vias_gen$8$2$2$1$2
X$10 VDD VDD \$25 OUT pfet$5$2$2$1$2
X$11 VDD VDD \$28 OUT pfet$5$2$2$1$2
X$12 OUT vias_gen$8$2$2$1$2
X$13 OUT vias_gen$12$2$2$1$2
X$14 IN OUT VDD VDD pfet$4$2$2$1$2
X$15 IN VDD OUT VDD pfet$4$2$2$1$2
X$16 OUT vias_gen$13$2$2$1$2
X$17 IN VDD OUT VDD pfet$4$2$2$1$2
X$18 OUT vias_gen$13$2$2$1$2
X$19 IN OUT VDD VDD pfet$4$2$2$1$2
X$20 OUT vias_gen$16$2$2$1$2
X$21 OUT vias_gen$16$2$2$1$2
X$22 IN vias_gen$14$2$2$1$2
X$23 IN vias_gen$14$2$2$1$2
X$24 IN vias_gen$14$2$2$1$2
X$25 IN vias_gen$14$2$2$1$2
X$26 VDD vias_gen$17$2$2$1$2
X$27 VDD vias_gen$17$2$2$1$2
X$28 VDD vias_gen$15$2$2$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$2$1$2

.SUBCKT rovcel2_LVT$1$1$2$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$2$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$2$1$2
X$3 IN GND OUT nfet$4$1$2$1$2
X$4 GND vias_gen$17$1$1$2$1$2
X$5 GND vias_gen$15$1$1$2$1$2
X$6 GND vias_gen$17$1$1$2$1$2
X$7 IN OUT GND nfet$4$1$2$1$2
X$8 OUT vias_gen$12$1$1$2$1$2
X$9 OUT vias_gen$8$1$1$2$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$1$2$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$1$2$1$2
X$12 OUT vias_gen$8$1$1$2$1$2
X$13 OUT vias_gen$12$1$1$2$1$2
X$14 OUT vias_gen$16$1$1$2$1$2
X$15 OUT vias_gen$16$1$1$2$1$2
X$16 IN OUT VDD VDD pfet$4$1$1$2$1$2
X$17 OUT vias_gen$13$1$1$2$1$2
X$18 IN VDD OUT VDD pfet$4$1$1$2$1$2
X$19 OUT vias_gen$13$1$1$2$1$2
X$20 IN VDD OUT VDD pfet$4$1$1$2$1$2
X$21 IN OUT VDD VDD pfet$4$1$1$2$1$2
X$22 IN vias_gen$14$1$1$2$1$2
X$23 IN vias_gen$14$1$1$2$1$2
X$24 IN vias_gen$14$1$1$2$1$2
X$25 IN vias_gen$14$1$1$2$1$2
X$26 VDD vias_gen$17$1$1$2$1$2
X$27 VDD vias_gen$15$1$1$2$1$2
X$28 VDD vias_gen$17$1$1$2$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$2$1$2

.SUBCKT rovcel2_LVT$2$1$2$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$2$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$2$2
X$3 IN OUT GND nfet$5$1$2$2
X$4 IN GND OUT nfet$5$1$2$2
X$5 GND vias_gen$17$2$1$2$2
X$6 GND vias_gen$17$2$1$2$2
X$7 GND vias_gen$15$2$1$2$2
X$8 OUT vias_gen$12$2$1$2$2
X$9 OUT vias_gen$8$2$1$2$2
X$10 VDD VDD \$25 OUT pfet$5$2$1$2$2
X$11 VDD VDD \$28 OUT pfet$5$2$1$2$2
X$12 OUT vias_gen$8$2$1$2$2
X$13 OUT vias_gen$12$2$1$2$2
X$14 IN OUT VDD VDD pfet$4$2$1$2$2
X$15 IN VDD OUT VDD pfet$4$2$1$2$2
X$16 OUT vias_gen$13$2$1$2$2
X$17 IN VDD OUT VDD pfet$4$2$1$2$2
X$18 OUT vias_gen$13$2$1$2$2
X$19 IN OUT VDD VDD pfet$4$2$1$2$2
X$20 OUT vias_gen$16$2$1$2$2
X$21 OUT vias_gen$16$2$1$2$2
X$22 IN vias_gen$14$2$1$2$2
X$23 IN vias_gen$14$2$1$2$2
X$24 IN vias_gen$14$2$1$2$2
X$25 IN vias_gen$14$2$1$2$2
X$26 VDD vias_gen$17$2$1$2$2
X$27 VDD vias_gen$17$2$1$2$2
X$28 VDD vias_gen$15$2$1$2$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$2$2

.SUBCKT rovcel2_LVT$1$1$1$2$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$2$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$2$2
X$3 IN GND OUT nfet$4$1$1$2$2
X$4 GND vias_gen$17$1$1$1$2$2
X$5 GND vias_gen$15$1$1$1$2$2
X$6 GND vias_gen$17$1$1$1$2$2
X$7 IN OUT GND nfet$4$1$1$2$2
X$8 OUT vias_gen$12$1$1$1$2$2
X$9 OUT vias_gen$8$1$1$1$2$2
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$2$2
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$2$2
X$12 OUT vias_gen$8$1$1$1$2$2
X$13 OUT vias_gen$12$1$1$1$2$2
X$14 OUT vias_gen$16$1$1$1$2$2
X$15 OUT vias_gen$16$1$1$1$2$2
X$16 IN OUT VDD VDD pfet$4$1$1$1$2$2
X$17 OUT vias_gen$13$1$1$1$2$2
X$18 IN VDD OUT VDD pfet$4$1$1$1$2$2
X$19 OUT vias_gen$13$1$1$1$2$2
X$20 IN VDD OUT VDD pfet$4$1$1$1$2$2
X$21 IN OUT VDD VDD pfet$4$1$1$1$2$2
X$22 IN vias_gen$14$1$1$1$2$2
X$23 IN vias_gen$14$1$1$1$2$2
X$24 IN vias_gen$14$1$1$1$2$2
X$25 IN vias_gen$14$1$1$1$2$2
X$26 VDD vias_gen$17$1$1$1$2$2
X$27 VDD vias_gen$15$1$1$1$2$2
X$28 VDD vias_gen$17$1$1$1$2$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$2$2

.SUBCKT rovcel2_LVT$3$2$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$2$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$2$2
X$3 IN OUT GND nfet$6$2$2
X$4 IN GND OUT nfet$6$2$2
X$5 GND vias_gen$17$3$2$2
X$6 GND vias_gen$17$3$2$2
X$7 GND vias_gen$15$3$2$2
X$8 OUT vias_gen$12$3$2$2
X$9 OUT vias_gen$8$3$2$2
X$10 VDD VDD \$25 OUT pfet$5$3$2$2
X$11 VDD VDD \$28 OUT pfet$5$3$2$2
X$12 OUT vias_gen$8$3$2$2
X$13 OUT vias_gen$12$3$2$2
X$14 IN OUT VDD VDD pfet$4$3$2$2
X$15 IN VDD OUT VDD pfet$4$3$2$2
X$16 OUT vias_gen$13$3$2$2
X$17 IN VDD OUT VDD pfet$4$3$2$2
X$18 OUT vias_gen$13$3$2$2
X$19 IN OUT VDD VDD pfet$4$3$2$2
X$20 OUT vias_gen$16$3$2$2
X$21 OUT vias_gen$16$3$2$2
X$22 IN vias_gen$14$3$2$2
X$23 IN vias_gen$14$3$2$2
X$24 IN vias_gen$14$3$2$2
X$25 IN vias_gen$14$3$2$2
X$26 VDD vias_gen$17$3$2$2
X$27 VDD vias_gen$17$3$2$2
X$28 VDD vias_gen$15$3$2$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$2$2

.SUBCKT rovcel2_LVT$1$2$2$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$2$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$2$2
X$3 IN GND OUT nfet$4$2$2$2
X$4 GND vias_gen$17$1$2$2$2
X$5 GND vias_gen$15$1$2$2$2
X$6 GND vias_gen$17$1$2$2$2
X$7 IN OUT GND nfet$4$2$2$2
X$8 OUT vias_gen$12$1$2$2$2
X$9 OUT vias_gen$8$1$2$2$2
X$10 VDD VDD \$25 OUT pfet$5$1$2$2$2
X$11 VDD VDD \$27 OUT pfet$5$1$2$2$2
X$12 OUT vias_gen$8$1$2$2$2
X$13 OUT vias_gen$12$1$2$2$2
X$14 OUT vias_gen$16$1$2$2$2
X$15 OUT vias_gen$16$1$2$2$2
X$16 IN OUT VDD VDD pfet$4$1$2$2$2
X$17 OUT vias_gen$13$1$2$2$2
X$18 IN VDD OUT VDD pfet$4$1$2$2$2
X$19 OUT vias_gen$13$1$2$2$2
X$20 IN VDD OUT VDD pfet$4$1$2$2$2
X$21 IN OUT VDD VDD pfet$4$1$2$2$2
X$22 IN vias_gen$14$1$2$2$2
X$23 IN vias_gen$14$1$2$2$2
X$24 IN vias_gen$14$1$2$2$2
X$25 IN vias_gen$14$1$2$2$2
X$26 VDD vias_gen$17$1$2$2$2
X$27 VDD vias_gen$15$1$2$2$2
X$28 VDD vias_gen$17$1$2$2$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$2$2

.SUBCKT rovcel2_LVT$3$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$1$1$1
X$3 IN OUT GND nfet$6$1$1$1
X$4 IN GND OUT nfet$6$1$1$1
X$5 GND vias_gen$17$3$1$1$1
X$6 GND vias_gen$17$3$1$1$1
X$7 GND vias_gen$15$3$1$1$1
X$8 OUT vias_gen$12$3$1$1$1
X$9 OUT vias_gen$8$3$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$3$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$3$1$1$1
X$12 OUT vias_gen$8$3$1$1$1
X$13 OUT vias_gen$12$3$1$1$1
X$14 IN OUT VDD VDD pfet$4$3$1$1$1
X$15 IN VDD OUT VDD pfet$4$3$1$1$1
X$16 OUT vias_gen$13$3$1$1$1
X$17 IN VDD OUT VDD pfet$4$3$1$1$1
X$18 OUT vias_gen$13$3$1$1$1
X$19 IN OUT VDD VDD pfet$4$3$1$1$1
X$20 OUT vias_gen$16$3$1$1$1
X$21 OUT vias_gen$16$3$1$1$1
X$22 IN vias_gen$14$3$1$1$1
X$23 IN vias_gen$14$3$1$1$1
X$24 IN vias_gen$14$3$1$1$1
X$25 IN vias_gen$14$3$1$1$1
X$26 VDD vias_gen$17$3$1$1$1
X$27 VDD vias_gen$17$3$1$1$1
X$28 VDD vias_gen$15$3$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$1$1$1

.SUBCKT rovcel2_LVT$1$2$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$1$1$1
X$3 IN GND OUT nfet$4$2$1$1$1
X$4 GND vias_gen$17$1$2$1$1$1
X$5 GND vias_gen$15$1$2$1$1$1
X$6 GND vias_gen$17$1$2$1$1$1
X$7 IN OUT GND nfet$4$2$1$1$1
X$8 OUT vias_gen$12$1$2$1$1$1
X$9 OUT vias_gen$8$1$2$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$2$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$2$1$1$1
X$12 OUT vias_gen$8$1$2$1$1$1
X$13 OUT vias_gen$12$1$2$1$1$1
X$14 OUT vias_gen$16$1$2$1$1$1
X$15 OUT vias_gen$16$1$2$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$2$1$1$1
X$17 OUT vias_gen$13$1$2$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$2$1$1$1
X$19 OUT vias_gen$13$1$2$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$2$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$2$1$1$1
X$22 IN vias_gen$14$1$2$1$1$1
X$23 IN vias_gen$14$1$2$1$1$1
X$24 IN vias_gen$14$1$2$1$1$1
X$25 IN vias_gen$14$1$2$1$1$1
X$26 VDD vias_gen$17$1$2$1$1$1
X$27 VDD vias_gen$15$1$2$1$1$1
X$28 VDD vias_gen$17$1$2$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$1$1$1

.SUBCKT rovcel2_LVT$2$2$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$2$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$2$1$1
X$3 IN OUT GND nfet$5$2$1$1
X$4 IN GND OUT nfet$5$2$1$1
X$5 GND vias_gen$17$2$2$1$1
X$6 GND vias_gen$17$2$2$1$1
X$7 GND vias_gen$15$2$2$1$1
X$8 OUT vias_gen$12$2$2$1$1
X$9 OUT vias_gen$8$2$2$1$1
X$10 VDD VDD \$25 OUT pfet$5$2$2$1$1
X$11 VDD VDD \$28 OUT pfet$5$2$2$1$1
X$12 OUT vias_gen$8$2$2$1$1
X$13 OUT vias_gen$12$2$2$1$1
X$14 IN OUT VDD VDD pfet$4$2$2$1$1
X$15 IN VDD OUT VDD pfet$4$2$2$1$1
X$16 OUT vias_gen$13$2$2$1$1
X$17 IN VDD OUT VDD pfet$4$2$2$1$1
X$18 OUT vias_gen$13$2$2$1$1
X$19 IN OUT VDD VDD pfet$4$2$2$1$1
X$20 OUT vias_gen$16$2$2$1$1
X$21 OUT vias_gen$16$2$2$1$1
X$22 IN vias_gen$14$2$2$1$1
X$23 IN vias_gen$14$2$2$1$1
X$24 IN vias_gen$14$2$2$1$1
X$25 IN vias_gen$14$2$2$1$1
X$26 VDD vias_gen$17$2$2$1$1
X$27 VDD vias_gen$17$2$2$1$1
X$28 VDD vias_gen$15$2$2$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$2$1$1

.SUBCKT rovcel2_LVT$1$1$2$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$2$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$2$1$1
X$3 IN GND OUT nfet$4$1$2$1$1
X$4 GND vias_gen$17$1$1$2$1$1
X$5 GND vias_gen$15$1$1$2$1$1
X$6 GND vias_gen$17$1$1$2$1$1
X$7 IN OUT GND nfet$4$1$2$1$1
X$8 OUT vias_gen$12$1$1$2$1$1
X$9 OUT vias_gen$8$1$1$2$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$2$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$2$1$1
X$12 OUT vias_gen$8$1$1$2$1$1
X$13 OUT vias_gen$12$1$1$2$1$1
X$14 OUT vias_gen$16$1$1$2$1$1
X$15 OUT vias_gen$16$1$1$2$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$2$1$1
X$17 OUT vias_gen$13$1$1$2$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$2$1$1
X$19 OUT vias_gen$13$1$1$2$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$2$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$2$1$1
X$22 IN vias_gen$14$1$1$2$1$1
X$23 IN vias_gen$14$1$1$2$1$1
X$24 IN vias_gen$14$1$1$2$1$1
X$25 IN vias_gen$14$1$1$2$1$1
X$26 VDD vias_gen$17$1$1$2$1$1
X$27 VDD vias_gen$15$1$1$2$1$1
X$28 VDD vias_gen$17$1$1$2$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$2$1$1

.SUBCKT rovcel2_LVT$2$1$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$2$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$2$1
X$3 IN OUT GND nfet$5$1$2$1
X$4 IN GND OUT nfet$5$1$2$1
X$5 GND vias_gen$17$2$1$2$1
X$6 GND vias_gen$17$2$1$2$1
X$7 GND vias_gen$15$2$1$2$1
X$8 OUT vias_gen$12$2$1$2$1
X$9 OUT vias_gen$8$2$1$2$1
X$10 VDD VDD \$25 OUT pfet$5$2$1$2$1
X$11 VDD VDD \$28 OUT pfet$5$2$1$2$1
X$12 OUT vias_gen$8$2$1$2$1
X$13 OUT vias_gen$12$2$1$2$1
X$14 IN OUT VDD VDD pfet$4$2$1$2$1
X$15 IN VDD OUT VDD pfet$4$2$1$2$1
X$16 OUT vias_gen$13$2$1$2$1
X$17 IN VDD OUT VDD pfet$4$2$1$2$1
X$18 OUT vias_gen$13$2$1$2$1
X$19 IN OUT VDD VDD pfet$4$2$1$2$1
X$20 OUT vias_gen$16$2$1$2$1
X$21 OUT vias_gen$16$2$1$2$1
X$22 IN vias_gen$14$2$1$2$1
X$23 IN vias_gen$14$2$1$2$1
X$24 IN vias_gen$14$2$1$2$1
X$25 IN vias_gen$14$2$1$2$1
X$26 VDD vias_gen$17$2$1$2$1
X$27 VDD vias_gen$17$2$1$2$1
X$28 VDD vias_gen$15$2$1$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$2$1

.SUBCKT rovcel2_LVT$1$1$1$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$2$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$2$1
X$3 IN GND OUT nfet$4$1$1$2$1
X$4 GND vias_gen$17$1$1$1$2$1
X$5 GND vias_gen$15$1$1$1$2$1
X$6 GND vias_gen$17$1$1$1$2$1
X$7 IN OUT GND nfet$4$1$1$2$1
X$8 OUT vias_gen$12$1$1$1$2$1
X$9 OUT vias_gen$8$1$1$1$2$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$2$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$2$1
X$12 OUT vias_gen$8$1$1$1$2$1
X$13 OUT vias_gen$12$1$1$1$2$1
X$14 OUT vias_gen$16$1$1$1$2$1
X$15 OUT vias_gen$16$1$1$1$2$1
X$16 IN OUT VDD VDD pfet$4$1$1$1$2$1
X$17 OUT vias_gen$13$1$1$1$2$1
X$18 IN VDD OUT VDD pfet$4$1$1$1$2$1
X$19 OUT vias_gen$13$1$1$1$2$1
X$20 IN VDD OUT VDD pfet$4$1$1$1$2$1
X$21 IN OUT VDD VDD pfet$4$1$1$1$2$1
X$22 IN vias_gen$14$1$1$1$2$1
X$23 IN vias_gen$14$1$1$1$2$1
X$24 IN vias_gen$14$1$1$1$2$1
X$25 IN vias_gen$14$1$1$1$2$1
X$26 VDD vias_gen$17$1$1$1$2$1
X$27 VDD vias_gen$15$1$1$1$2$1
X$28 VDD vias_gen$17$1$1$1$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$2$1

.SUBCKT rovcel2_LVT$3$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$2$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$2$1
X$3 IN OUT GND nfet$6$2$1
X$4 IN GND OUT nfet$6$2$1
X$5 GND vias_gen$17$3$2$1
X$6 GND vias_gen$17$3$2$1
X$7 GND vias_gen$15$3$2$1
X$8 OUT vias_gen$12$3$2$1
X$9 OUT vias_gen$8$3$2$1
X$10 VDD VDD \$25 OUT pfet$5$3$2$1
X$11 VDD VDD \$28 OUT pfet$5$3$2$1
X$12 OUT vias_gen$8$3$2$1
X$13 OUT vias_gen$12$3$2$1
X$14 IN OUT VDD VDD pfet$4$3$2$1
X$15 IN VDD OUT VDD pfet$4$3$2$1
X$16 OUT vias_gen$13$3$2$1
X$17 IN VDD OUT VDD pfet$4$3$2$1
X$18 OUT vias_gen$13$3$2$1
X$19 IN OUT VDD VDD pfet$4$3$2$1
X$20 OUT vias_gen$16$3$2$1
X$21 OUT vias_gen$16$3$2$1
X$22 IN vias_gen$14$3$2$1
X$23 IN vias_gen$14$3$2$1
X$24 IN vias_gen$14$3$2$1
X$25 IN vias_gen$14$3$2$1
X$26 VDD vias_gen$17$3$2$1
X$27 VDD vias_gen$17$3$2$1
X$28 VDD vias_gen$15$3$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$2$1

.SUBCKT rovcel2_LVT$1$2$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$2$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$2$1
X$3 IN GND OUT nfet$4$2$2$1
X$4 GND vias_gen$17$1$2$2$1
X$5 GND vias_gen$15$1$2$2$1
X$6 GND vias_gen$17$1$2$2$1
X$7 IN OUT GND nfet$4$2$2$1
X$8 OUT vias_gen$12$1$2$2$1
X$9 OUT vias_gen$8$1$2$2$1
X$10 VDD VDD \$25 OUT pfet$5$1$2$2$1
X$11 VDD VDD \$27 OUT pfet$5$1$2$2$1
X$12 OUT vias_gen$8$1$2$2$1
X$13 OUT vias_gen$12$1$2$2$1
X$14 OUT vias_gen$16$1$2$2$1
X$15 OUT vias_gen$16$1$2$2$1
X$16 IN OUT VDD VDD pfet$4$1$2$2$1
X$17 OUT vias_gen$13$1$2$2$1
X$18 IN VDD OUT VDD pfet$4$1$2$2$1
X$19 OUT vias_gen$13$1$2$2$1
X$20 IN VDD OUT VDD pfet$4$1$2$2$1
X$21 IN OUT VDD VDD pfet$4$1$2$2$1
X$22 IN vias_gen$14$1$2$2$1
X$23 IN vias_gen$14$1$2$2$1
X$24 IN vias_gen$14$1$2$2$1
X$25 IN vias_gen$14$1$2$2$1
X$26 VDD vias_gen$17$1$2$2$1
X$27 VDD vias_gen$15$1$2$2$1
X$28 VDD vias_gen$17$1$2$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$2$1

.SUBCKT rovcel2_LVT$2$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$1$1
X$3 IN OUT GND nfet$5$1$1$1
X$4 IN GND OUT nfet$5$1$1$1
X$5 GND vias_gen$17$2$1$1$1
X$6 GND vias_gen$17$2$1$1$1
X$7 GND vias_gen$15$2$1$1$1
X$8 OUT vias_gen$12$2$1$1$1
X$9 OUT vias_gen$8$2$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$2$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$2$1$1$1
X$12 OUT vias_gen$8$2$1$1$1
X$13 OUT vias_gen$12$2$1$1$1
X$14 IN OUT VDD VDD pfet$4$2$1$1$1
X$15 IN VDD OUT VDD pfet$4$2$1$1$1
X$16 OUT vias_gen$13$2$1$1$1
X$17 IN VDD OUT VDD pfet$4$2$1$1$1
X$18 OUT vias_gen$13$2$1$1$1
X$19 IN OUT VDD VDD pfet$4$2$1$1$1
X$20 OUT vias_gen$16$2$1$1$1
X$21 OUT vias_gen$16$2$1$1$1
X$22 IN vias_gen$14$2$1$1$1
X$23 IN vias_gen$14$2$1$1$1
X$24 IN vias_gen$14$2$1$1$1
X$25 IN vias_gen$14$2$1$1$1
X$26 VDD vias_gen$17$2$1$1$1
X$27 VDD vias_gen$17$2$1$1$1
X$28 VDD vias_gen$15$2$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$1$1

.SUBCKT rovcel2_LVT$1$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$1$1
X$3 IN GND OUT nfet$4$1$1$1$1
X$4 GND vias_gen$17$1$1$1$1$1
X$5 GND vias_gen$15$1$1$1$1$1
X$6 GND vias_gen$17$1$1$1$1$1
X$7 IN OUT GND nfet$4$1$1$1$1
X$8 OUT vias_gen$12$1$1$1$1$1
X$9 OUT vias_gen$8$1$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$1$1
X$12 OUT vias_gen$8$1$1$1$1$1
X$13 OUT vias_gen$12$1$1$1$1$1
X$14 OUT vias_gen$16$1$1$1$1$1
X$15 OUT vias_gen$16$1$1$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$1$1$1
X$17 OUT vias_gen$13$1$1$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$1$1$1
X$19 OUT vias_gen$13$1$1$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$1$1$1
X$22 IN vias_gen$14$1$1$1$1$1
X$23 IN vias_gen$14$1$1$1$1$1
X$24 IN vias_gen$14$1$1$1$1$1
X$25 IN vias_gen$14$1$1$1$1$1
X$26 VDD vias_gen$17$1$1$1$1$1
X$27 VDD vias_gen$15$1$1$1$1$1
X$28 VDD vias_gen$17$1$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$1$1

.SUBCKT rovcel2_LVT$3$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$1$1
X$3 IN OUT GND nfet$6$1$1
X$4 IN GND OUT nfet$6$1$1
X$5 GND vias_gen$17$3$1$1
X$6 GND vias_gen$17$3$1$1
X$7 GND vias_gen$15$3$1$1
X$8 OUT vias_gen$12$3$1$1
X$9 OUT vias_gen$8$3$1$1
X$10 VDD VDD \$25 OUT pfet$5$3$1$1
X$11 VDD VDD \$28 OUT pfet$5$3$1$1
X$12 OUT vias_gen$8$3$1$1
X$13 OUT vias_gen$12$3$1$1
X$14 IN OUT VDD VDD pfet$4$3$1$1
X$15 IN VDD OUT VDD pfet$4$3$1$1
X$16 OUT vias_gen$13$3$1$1
X$17 IN VDD OUT VDD pfet$4$3$1$1
X$18 OUT vias_gen$13$3$1$1
X$19 IN OUT VDD VDD pfet$4$3$1$1
X$20 OUT vias_gen$16$3$1$1
X$21 OUT vias_gen$16$3$1$1
X$22 IN vias_gen$14$3$1$1
X$23 IN vias_gen$14$3$1$1
X$24 IN vias_gen$14$3$1$1
X$25 IN vias_gen$14$3$1$1
X$26 VDD vias_gen$17$3$1$1
X$27 VDD vias_gen$17$3$1$1
X$28 VDD vias_gen$15$3$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$1$1

.SUBCKT rovcel2_LVT$1$2$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$1$1
X$3 IN GND OUT nfet$4$2$1$1
X$4 GND vias_gen$17$1$2$1$1
X$5 GND vias_gen$15$1$2$1$1
X$6 GND vias_gen$17$1$2$1$1
X$7 IN OUT GND nfet$4$2$1$1
X$8 OUT vias_gen$12$1$2$1$1
X$9 OUT vias_gen$8$1$2$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$2$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$2$1$1
X$12 OUT vias_gen$8$1$2$1$1
X$13 OUT vias_gen$12$1$2$1$1
X$14 OUT vias_gen$16$1$2$1$1
X$15 OUT vias_gen$16$1$2$1$1
X$16 IN OUT VDD VDD pfet$4$1$2$1$1
X$17 OUT vias_gen$13$1$2$1$1
X$18 IN VDD OUT VDD pfet$4$1$2$1$1
X$19 OUT vias_gen$13$1$2$1$1
X$20 IN VDD OUT VDD pfet$4$1$2$1$1
X$21 IN OUT VDD VDD pfet$4$1$2$1$1
X$22 IN vias_gen$14$1$2$1$1
X$23 IN vias_gen$14$1$2$1$1
X$24 IN vias_gen$14$1$2$1$1
X$25 IN vias_gen$14$1$2$1$1
X$26 VDD vias_gen$17$1$2$1$1
X$27 VDD vias_gen$15$1$2$1$1
X$28 VDD vias_gen$17$1$2$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$1$1

.SUBCKT rovcel2_LVT$2$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$2$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$2$1
X$3 IN OUT GND nfet$5$2$1
X$4 IN GND OUT nfet$5$2$1
X$5 GND vias_gen$17$2$2$1
X$6 GND vias_gen$17$2$2$1
X$7 GND vias_gen$15$2$2$1
X$8 OUT vias_gen$12$2$2$1
X$9 OUT vias_gen$8$2$2$1
X$10 VDD VDD \$25 OUT pfet$5$2$2$1
X$11 VDD VDD \$28 OUT pfet$5$2$2$1
X$12 OUT vias_gen$8$2$2$1
X$13 OUT vias_gen$12$2$2$1
X$14 IN OUT VDD VDD pfet$4$2$2$1
X$15 IN VDD OUT VDD pfet$4$2$2$1
X$16 OUT vias_gen$13$2$2$1
X$17 IN VDD OUT VDD pfet$4$2$2$1
X$18 OUT vias_gen$13$2$2$1
X$19 IN OUT VDD VDD pfet$4$2$2$1
X$20 OUT vias_gen$16$2$2$1
X$21 OUT vias_gen$16$2$2$1
X$22 IN vias_gen$14$2$2$1
X$23 IN vias_gen$14$2$2$1
X$24 IN vias_gen$14$2$2$1
X$25 IN vias_gen$14$2$2$1
X$26 VDD vias_gen$17$2$2$1
X$27 VDD vias_gen$17$2$2$1
X$28 VDD vias_gen$15$2$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$2$1

.SUBCKT rovcel2_LVT$1$1$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$2$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$2$1
X$3 IN GND OUT nfet$4$1$2$1
X$4 GND vias_gen$17$1$1$2$1
X$5 GND vias_gen$15$1$1$2$1
X$6 GND vias_gen$17$1$1$2$1
X$7 IN OUT GND nfet$4$1$2$1
X$8 OUT vias_gen$12$1$1$2$1
X$9 OUT vias_gen$8$1$1$2$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$2$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$2$1
X$12 OUT vias_gen$8$1$1$2$1
X$13 OUT vias_gen$12$1$1$2$1
X$14 OUT vias_gen$16$1$1$2$1
X$15 OUT vias_gen$16$1$1$2$1
X$16 IN OUT VDD VDD pfet$4$1$1$2$1
X$17 OUT vias_gen$13$1$1$2$1
X$18 IN VDD OUT VDD pfet$4$1$1$2$1
X$19 OUT vias_gen$13$1$1$2$1
X$20 IN VDD OUT VDD pfet$4$1$1$2$1
X$21 IN OUT VDD VDD pfet$4$1$1$2$1
X$22 IN vias_gen$14$1$1$2$1
X$23 IN vias_gen$14$1$1$2$1
X$24 IN vias_gen$14$1$1$2$1
X$25 IN vias_gen$14$1$1$2$1
X$26 VDD vias_gen$17$1$1$2$1
X$27 VDD vias_gen$15$1$1$2$1
X$28 VDD vias_gen$17$1$1$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$2$1

.SUBCKT rovcel2_LVT$2$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$2
X$3 IN OUT GND nfet$5$1$2
X$4 IN GND OUT nfet$5$1$2
X$5 GND vias_gen$17$2$1$2
X$6 GND vias_gen$17$2$1$2
X$7 GND vias_gen$15$2$1$2
X$8 OUT vias_gen$12$2$1$2
X$9 OUT vias_gen$8$2$1$2
X$10 VDD VDD \$25 OUT pfet$5$2$1$2
X$11 VDD VDD \$28 OUT pfet$5$2$1$2
X$12 OUT vias_gen$8$2$1$2
X$13 OUT vias_gen$12$2$1$2
X$14 IN OUT VDD VDD pfet$4$2$1$2
X$15 IN VDD OUT VDD pfet$4$2$1$2
X$16 OUT vias_gen$13$2$1$2
X$17 IN VDD OUT VDD pfet$4$2$1$2
X$18 OUT vias_gen$13$2$1$2
X$19 IN OUT VDD VDD pfet$4$2$1$2
X$20 OUT vias_gen$16$2$1$2
X$21 OUT vias_gen$16$2$1$2
X$22 IN vias_gen$14$2$1$2
X$23 IN vias_gen$14$2$1$2
X$24 IN vias_gen$14$2$1$2
X$25 IN vias_gen$14$2$1$2
X$26 VDD vias_gen$17$2$1$2
X$27 VDD vias_gen$17$2$1$2
X$28 VDD vias_gen$15$2$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$2

.SUBCKT rovcel2_LVT$1$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$2
X$3 IN GND OUT nfet$4$1$1$2
X$4 GND vias_gen$17$1$1$1$2
X$5 GND vias_gen$15$1$1$1$2
X$6 GND vias_gen$17$1$1$1$2
X$7 IN OUT GND nfet$4$1$1$2
X$8 OUT vias_gen$12$1$1$1$2
X$9 OUT vias_gen$8$1$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$2
X$12 OUT vias_gen$8$1$1$1$2
X$13 OUT vias_gen$12$1$1$1$2
X$14 OUT vias_gen$16$1$1$1$2
X$15 OUT vias_gen$16$1$1$1$2
X$16 IN OUT VDD VDD pfet$4$1$1$1$2
X$17 OUT vias_gen$13$1$1$1$2
X$18 IN VDD OUT VDD pfet$4$1$1$1$2
X$19 OUT vias_gen$13$1$1$1$2
X$20 IN VDD OUT VDD pfet$4$1$1$1$2
X$21 IN OUT VDD VDD pfet$4$1$1$1$2
X$22 IN vias_gen$14$1$1$1$2
X$23 IN vias_gen$14$1$1$1$2
X$24 IN vias_gen$14$1$1$1$2
X$25 IN vias_gen$14$1$1$1$2
X$26 VDD vias_gen$17$1$1$1$2
X$27 VDD vias_gen$15$1$1$1$2
X$28 VDD vias_gen$17$1$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$2

.SUBCKT rovcel2_LVT$3$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$2
X$3 IN OUT GND nfet$6$2
X$4 IN GND OUT nfet$6$2
X$5 GND vias_gen$17$3$2
X$6 GND vias_gen$17$3$2
X$7 GND vias_gen$15$3$2
X$8 OUT vias_gen$12$3$2
X$9 OUT vias_gen$8$3$2
X$10 VDD VDD \$25 OUT pfet$5$3$2
X$11 VDD VDD \$28 OUT pfet$5$3$2
X$12 OUT vias_gen$8$3$2
X$13 OUT vias_gen$12$3$2
X$14 IN OUT VDD VDD pfet$4$3$2
X$15 IN VDD OUT VDD pfet$4$3$2
X$16 OUT vias_gen$13$3$2
X$17 IN VDD OUT VDD pfet$4$3$2
X$18 OUT vias_gen$13$3$2
X$19 IN OUT VDD VDD pfet$4$3$2
X$20 OUT vias_gen$16$3$2
X$21 OUT vias_gen$16$3$2
X$22 IN vias_gen$14$3$2
X$23 IN vias_gen$14$3$2
X$24 IN vias_gen$14$3$2
X$25 IN vias_gen$14$3$2
X$26 VDD vias_gen$17$3$2
X$27 VDD vias_gen$17$3$2
X$28 VDD vias_gen$15$3$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$2

.SUBCKT rovcel2_LVT$1$2$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$2
X$3 IN GND OUT nfet$4$2$2
X$4 GND vias_gen$17$1$2$2
X$5 GND vias_gen$15$1$2$2
X$6 GND vias_gen$17$1$2$2
X$7 IN OUT GND nfet$4$2$2
X$8 OUT vias_gen$12$1$2$2
X$9 OUT vias_gen$8$1$2$2
X$10 VDD VDD \$25 OUT pfet$5$1$2$2
X$11 VDD VDD \$27 OUT pfet$5$1$2$2
X$12 OUT vias_gen$8$1$2$2
X$13 OUT vias_gen$12$1$2$2
X$14 OUT vias_gen$16$1$2$2
X$15 OUT vias_gen$16$1$2$2
X$16 IN OUT VDD VDD pfet$4$1$2$2
X$17 OUT vias_gen$13$1$2$2
X$18 IN VDD OUT VDD pfet$4$1$2$2
X$19 OUT vias_gen$13$1$2$2
X$20 IN VDD OUT VDD pfet$4$1$2$2
X$21 IN OUT VDD VDD pfet$4$1$2$2
X$22 IN vias_gen$14$1$2$2
X$23 IN vias_gen$14$1$2$2
X$24 IN vias_gen$14$1$2$2
X$25 IN vias_gen$14$1$2$2
X$26 VDD vias_gen$17$1$2$2
X$27 VDD vias_gen$15$1$2$2
X$28 VDD vias_gen$17$1$2$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$2

.SUBCKT rovcel2_LVT$2$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$1
X$3 IN OUT GND nfet$5$1$1
X$4 IN GND OUT nfet$5$1$1
X$5 GND vias_gen$17$2$1$1
X$6 GND vias_gen$17$2$1$1
X$7 GND vias_gen$15$2$1$1
X$8 OUT vias_gen$12$2$1$1
X$9 OUT vias_gen$8$2$1$1
X$10 VDD VDD \$25 OUT pfet$5$2$1$1
X$11 VDD VDD \$28 OUT pfet$5$2$1$1
X$12 OUT vias_gen$8$2$1$1
X$13 OUT vias_gen$12$2$1$1
X$14 IN OUT VDD VDD pfet$4$2$1$1
X$15 IN VDD OUT VDD pfet$4$2$1$1
X$16 OUT vias_gen$13$2$1$1
X$17 IN VDD OUT VDD pfet$4$2$1$1
X$18 OUT vias_gen$13$2$1$1
X$19 IN OUT VDD VDD pfet$4$2$1$1
X$20 OUT vias_gen$16$2$1$1
X$21 OUT vias_gen$16$2$1$1
X$22 IN vias_gen$14$2$1$1
X$23 IN vias_gen$14$2$1$1
X$24 IN vias_gen$14$2$1$1
X$25 IN vias_gen$14$2$1$1
X$26 VDD vias_gen$17$2$1$1
X$27 VDD vias_gen$17$2$1$1
X$28 VDD vias_gen$15$2$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$1

.SUBCKT rovcel2_LVT$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$1
X$3 IN GND OUT nfet$4$1$1$1
X$4 GND vias_gen$17$1$1$1$1
X$5 GND vias_gen$15$1$1$1$1
X$6 GND vias_gen$17$1$1$1$1
X$7 IN OUT GND nfet$4$1$1$1
X$8 OUT vias_gen$12$1$1$1$1
X$9 OUT vias_gen$8$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$1
X$12 OUT vias_gen$8$1$1$1$1
X$13 OUT vias_gen$12$1$1$1$1
X$14 OUT vias_gen$16$1$1$1$1
X$15 OUT vias_gen$16$1$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$1$1
X$17 OUT vias_gen$13$1$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$1$1
X$19 OUT vias_gen$13$1$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$1$1
X$22 IN vias_gen$14$1$1$1$1
X$23 IN vias_gen$14$1$1$1$1
X$24 IN vias_gen$14$1$1$1$1
X$25 IN vias_gen$14$1$1$1$1
X$26 VDD vias_gen$17$1$1$1$1
X$27 VDD vias_gen$15$1$1$1$1
X$28 VDD vias_gen$17$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$1

.SUBCKT rovcel2_LVT$3$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3$1
X$3 IN OUT GND nfet$6$1
X$4 IN GND OUT nfet$6$1
X$5 GND vias_gen$17$3$1
X$6 GND vias_gen$17$3$1
X$7 GND vias_gen$15$3$1
X$8 OUT vias_gen$12$3$1
X$9 OUT vias_gen$8$3$1
X$10 VDD VDD \$25 OUT pfet$5$3$1
X$11 VDD VDD \$28 OUT pfet$5$3$1
X$12 OUT vias_gen$8$3$1
X$13 OUT vias_gen$12$3$1
X$14 IN OUT VDD VDD pfet$4$3$1
X$15 IN VDD OUT VDD pfet$4$3$1
X$16 OUT vias_gen$13$3$1
X$17 IN VDD OUT VDD pfet$4$3$1
X$18 OUT vias_gen$13$3$1
X$19 IN OUT VDD VDD pfet$4$3$1
X$20 OUT vias_gen$16$3$1
X$21 OUT vias_gen$16$3$1
X$22 IN vias_gen$14$3$1
X$23 IN vias_gen$14$3$1
X$24 IN vias_gen$14$3$1
X$25 IN vias_gen$14$3$1
X$26 VDD vias_gen$17$3$1
X$27 VDD vias_gen$17$3$1
X$28 VDD vias_gen$15$3$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3$1

.SUBCKT rovcel2_LVT$1$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2$1
X$3 IN GND OUT nfet$4$2$1
X$4 GND vias_gen$17$1$2$1
X$5 GND vias_gen$15$1$2$1
X$6 GND vias_gen$17$1$2$1
X$7 IN OUT GND nfet$4$2$1
X$8 OUT vias_gen$12$1$2$1
X$9 OUT vias_gen$8$1$2$1
X$10 VDD VDD \$25 OUT pfet$5$1$2$1
X$11 VDD VDD \$27 OUT pfet$5$1$2$1
X$12 OUT vias_gen$8$1$2$1
X$13 OUT vias_gen$12$1$2$1
X$14 OUT vias_gen$16$1$2$1
X$15 OUT vias_gen$16$1$2$1
X$16 IN OUT VDD VDD pfet$4$1$2$1
X$17 OUT vias_gen$13$1$2$1
X$18 IN VDD OUT VDD pfet$4$1$2$1
X$19 OUT vias_gen$13$1$2$1
X$20 IN VDD OUT VDD pfet$4$1$2$1
X$21 IN OUT VDD VDD pfet$4$1$2$1
X$22 IN vias_gen$14$1$2$1
X$23 IN vias_gen$14$1$2$1
X$24 IN vias_gen$14$1$2$1
X$25 IN vias_gen$14$1$2$1
X$26 VDD vias_gen$17$1$2$1
X$27 VDD vias_gen$15$1$2$1
X$28 VDD vias_gen$17$1$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2$1

.SUBCKT rovcel2_LVT$2$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$2
X$3 IN OUT GND nfet$5$2
X$4 IN GND OUT nfet$5$2
X$5 GND vias_gen$17$2$2
X$6 GND vias_gen$17$2$2
X$7 GND vias_gen$15$2$2
X$8 OUT vias_gen$12$2$2
X$9 OUT vias_gen$8$2$2
X$10 VDD VDD \$25 OUT pfet$5$2$2
X$11 VDD VDD \$28 OUT pfet$5$2$2
X$12 OUT vias_gen$8$2$2
X$13 OUT vias_gen$12$2$2
X$14 IN OUT VDD VDD pfet$4$2$2
X$15 IN VDD OUT VDD pfet$4$2$2
X$16 OUT vias_gen$13$2$2
X$17 IN VDD OUT VDD pfet$4$2$2
X$18 OUT vias_gen$13$2$2
X$19 IN OUT VDD VDD pfet$4$2$2
X$20 OUT vias_gen$16$2$2
X$21 OUT vias_gen$16$2$2
X$22 IN vias_gen$14$2$2
X$23 IN vias_gen$14$2$2
X$24 IN vias_gen$14$2$2
X$25 IN vias_gen$14$2$2
X$26 VDD vias_gen$17$2$2
X$27 VDD vias_gen$17$2$2
X$28 VDD vias_gen$15$2$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$2

.SUBCKT rovcel2_LVT$1$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$2
X$3 IN GND OUT nfet$4$1$2
X$4 GND vias_gen$17$1$1$2
X$5 GND vias_gen$15$1$1$2
X$6 GND vias_gen$17$1$1$2
X$7 IN OUT GND nfet$4$1$2
X$8 OUT vias_gen$12$1$1$2
X$9 OUT vias_gen$8$1$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$1$2
X$12 OUT vias_gen$8$1$1$2
X$13 OUT vias_gen$12$1$1$2
X$14 OUT vias_gen$16$1$1$2
X$15 OUT vias_gen$16$1$1$2
X$16 IN OUT VDD VDD pfet$4$1$1$2
X$17 OUT vias_gen$13$1$1$2
X$18 IN VDD OUT VDD pfet$4$1$1$2
X$19 OUT vias_gen$13$1$1$2
X$20 IN VDD OUT VDD pfet$4$1$1$2
X$21 IN OUT VDD VDD pfet$4$1$1$2
X$22 IN vias_gen$14$1$1$2
X$23 IN vias_gen$14$1$1$2
X$24 IN vias_gen$14$1$1$2
X$25 IN vias_gen$14$1$1$2
X$26 VDD vias_gen$17$1$1$2
X$27 VDD vias_gen$15$1$1$2
X$28 VDD vias_gen$17$1$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$2

.SUBCKT rovcel2_LVT$2$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1
X$3 IN OUT GND nfet$5$1
X$4 IN GND OUT nfet$5$1
X$5 GND vias_gen$17$2$1
X$6 GND vias_gen$17$2$1
X$7 GND vias_gen$15$2$1
X$8 OUT vias_gen$12$2$1
X$9 OUT vias_gen$8$2$1
X$10 VDD VDD \$25 OUT pfet$5$2$1
X$11 VDD VDD \$28 OUT pfet$5$2$1
X$12 OUT vias_gen$8$2$1
X$13 OUT vias_gen$12$2$1
X$14 IN OUT VDD VDD pfet$4$2$1
X$15 IN VDD OUT VDD pfet$4$2$1
X$16 OUT vias_gen$13$2$1
X$17 IN VDD OUT VDD pfet$4$2$1
X$18 OUT vias_gen$13$2$1
X$19 IN OUT VDD VDD pfet$4$2$1
X$20 OUT vias_gen$16$2$1
X$21 OUT vias_gen$16$2$1
X$22 IN vias_gen$14$2$1
X$23 IN vias_gen$14$2$1
X$24 IN vias_gen$14$2$1
X$25 IN vias_gen$14$2$1
X$26 VDD vias_gen$17$2$1
X$27 VDD vias_gen$17$2$1
X$28 VDD vias_gen$15$2$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1

.SUBCKT rovcel2_LVT$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1
X$3 IN GND OUT nfet$4$1$1
X$4 GND vias_gen$17$1$1$1
X$5 GND vias_gen$15$1$1$1
X$6 GND vias_gen$17$1$1$1
X$7 IN OUT GND nfet$4$1$1
X$8 OUT vias_gen$12$1$1$1
X$9 OUT vias_gen$8$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1
X$12 OUT vias_gen$8$1$1$1
X$13 OUT vias_gen$12$1$1$1
X$14 OUT vias_gen$16$1$1$1
X$15 OUT vias_gen$16$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$1
X$17 OUT vias_gen$13$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$1
X$19 OUT vias_gen$13$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$1
X$22 IN vias_gen$14$1$1$1
X$23 IN vias_gen$14$1$1$1
X$24 IN vias_gen$14$1$1$1
X$25 IN vias_gen$14$1$1$1
X$26 VDD vias_gen$17$1$1$1
X$27 VDD vias_gen$15$1$1$1
X$28 VDD vias_gen$17$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1

.SUBCKT rovcel2_LVT$3 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$3
X$2 GND GND \$28 OUT sky130_gnd nfet$3$3
X$3 IN OUT GND nfet$6
X$4 IN GND OUT nfet$6
X$5 GND vias_gen$17$3
X$6 GND vias_gen$17$3
X$7 GND vias_gen$15$3
X$8 OUT vias_gen$12$3
X$9 OUT vias_gen$8$3
X$10 VDD VDD \$25 OUT pfet$5$3
X$11 VDD VDD \$28 OUT pfet$5$3
X$12 OUT vias_gen$8$3
X$13 OUT vias_gen$12$3
X$14 IN OUT VDD VDD pfet$4$3
X$15 IN VDD OUT VDD pfet$4$3
X$16 OUT vias_gen$13$3
X$17 IN VDD OUT VDD pfet$4$3
X$18 OUT vias_gen$13$3
X$19 IN OUT VDD VDD pfet$4$3
X$20 OUT vias_gen$16$3
X$21 OUT vias_gen$16$3
X$22 IN vias_gen$14$3
X$23 IN vias_gen$14$3
X$24 IN vias_gen$14$3
X$25 IN vias_gen$14$3
X$26 VDD vias_gen$17$3
X$27 VDD vias_gen$17$3
X$28 VDD vias_gen$15$3
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$3

.SUBCKT rovcel2_LVT$1$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$2
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$2
X$3 IN GND OUT nfet$4$2
X$4 GND vias_gen$17$1$2
X$5 GND vias_gen$15$1$2
X$6 GND vias_gen$17$1$2
X$7 IN OUT GND nfet$4$2
X$8 OUT vias_gen$12$1$2
X$9 OUT vias_gen$8$1$2
X$10 VDD VDD \$25 OUT pfet$5$1$2
X$11 VDD VDD \$27 OUT pfet$5$1$2
X$12 OUT vias_gen$8$1$2
X$13 OUT vias_gen$12$1$2
X$14 OUT vias_gen$16$1$2
X$15 OUT vias_gen$16$1$2
X$16 IN OUT VDD VDD pfet$4$1$2
X$17 OUT vias_gen$13$1$2
X$18 IN VDD OUT VDD pfet$4$1$2
X$19 OUT vias_gen$13$1$2
X$20 IN VDD OUT VDD pfet$4$1$2
X$21 IN OUT VDD VDD pfet$4$1$2
X$22 IN vias_gen$14$1$2
X$23 IN vias_gen$14$1$2
X$24 IN vias_gen$14$1$2
X$25 IN vias_gen$14$1$2
X$26 VDD vias_gen$17$1$2
X$27 VDD vias_gen$15$1$2
X$28 VDD vias_gen$17$1$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$2

.SUBCKT rovcel2_LVT$2 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2
X$3 IN OUT GND nfet$5
X$4 IN GND OUT nfet$5
X$5 GND vias_gen$17$2
X$6 GND vias_gen$17$2
X$7 GND vias_gen$15$2
X$8 OUT vias_gen$12$2
X$9 OUT vias_gen$8$2
X$10 VDD VDD \$25 OUT pfet$5$2
X$11 VDD VDD \$28 OUT pfet$5$2
X$12 OUT vias_gen$8$2
X$13 OUT vias_gen$12$2
X$14 IN OUT VDD VDD pfet$4$2
X$15 IN VDD OUT VDD pfet$4$2
X$16 OUT vias_gen$13$2
X$17 IN VDD OUT VDD pfet$4$2
X$18 OUT vias_gen$13$2
X$19 IN OUT VDD VDD pfet$4$2
X$20 OUT vias_gen$16$2
X$21 OUT vias_gen$16$2
X$22 IN vias_gen$14$2
X$23 IN vias_gen$14$2
X$24 IN vias_gen$14$2
X$25 IN vias_gen$14$2
X$26 VDD vias_gen$17$2
X$27 VDD vias_gen$17$2
X$28 VDD vias_gen$15$2
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2

.SUBCKT rovcel2_LVT$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1
X$3 IN GND OUT nfet$4$1
X$4 GND vias_gen$17$1$1
X$5 GND vias_gen$15$1$1
X$6 GND vias_gen$17$1$1
X$7 IN OUT GND nfet$4$1
X$8 OUT vias_gen$12$1$1
X$9 OUT vias_gen$8$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1
X$12 OUT vias_gen$8$1$1
X$13 OUT vias_gen$12$1$1
X$14 OUT vias_gen$16$1$1
X$15 OUT vias_gen$16$1$1
X$16 IN OUT VDD VDD pfet$4$1$1
X$17 OUT vias_gen$13$1$1
X$18 IN VDD OUT VDD pfet$4$1$1
X$19 OUT vias_gen$13$1$1
X$20 IN VDD OUT VDD pfet$4$1$1
X$21 IN OUT VDD VDD pfet$4$1$1
X$22 IN vias_gen$14$1$1
X$23 IN vias_gen$14$1$1
X$24 IN vias_gen$14$1$1
X$25 IN vias_gen$14$1$1
X$26 VDD vias_gen$17$1$1
X$27 VDD vias_gen$15$1$1
X$28 VDD vias_gen$17$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1

.SUBCKT rovcel2_LVT GND IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3
X$2 GND GND \$28 OUT sky130_gnd nfet$3
X$3 IN OUT GND nfet
X$4 IN GND OUT nfet
X$5 GND vias_gen$17
X$6 GND vias_gen$17
X$7 GND vias_gen$15
X$8 OUT vias_gen$12
X$9 OUT vias_gen$8
X$10 VDD VDD \$25 OUT pfet$5
X$11 VDD VDD \$28 OUT pfet$5
X$12 OUT vias_gen$8
X$13 OUT vias_gen$12
X$14 IN OUT VDD VDD pfet$4
X$15 IN VDD OUT VDD pfet$4
X$16 OUT vias_gen$13
X$17 IN VDD OUT VDD pfet$4
X$18 OUT vias_gen$13
X$19 IN OUT VDD VDD pfet$4
X$20 OUT vias_gen$16
X$21 OUT vias_gen$16
X$22 IN vias_gen$14
X$23 IN vias_gen$14
X$24 IN vias_gen$14
X$25 IN vias_gen$14
X$26 VDD vias_gen$17
X$27 VDD vias_gen$17
X$28 VDD vias_gen$15
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT

.SUBCKT rovcel2_LVT$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1
X$3 IN GND OUT nfet$4
X$4 GND vias_gen$17$1
X$5 GND vias_gen$15$1
X$6 GND vias_gen$17$1
X$7 IN OUT GND nfet$4
X$8 OUT vias_gen$12$1
X$9 OUT vias_gen$8$1
X$10 VDD VDD \$25 OUT pfet$5$1
X$11 VDD VDD \$27 OUT pfet$5$1
X$12 OUT vias_gen$8$1
X$13 OUT vias_gen$12$1
X$14 OUT vias_gen$16$1
X$15 OUT vias_gen$16$1
X$16 IN OUT VDD VDD pfet$4$1
X$17 OUT vias_gen$13$1
X$18 IN VDD OUT VDD pfet$4$1
X$19 OUT vias_gen$13$1
X$20 IN VDD OUT VDD pfet$4$1
X$21 IN OUT VDD VDD pfet$4$1
X$22 IN vias_gen$14$1
X$23 IN vias_gen$14$1
X$24 IN vias_gen$14$1
X$25 IN vias_gen$14$1
X$26 VDD vias_gen$17$1
X$27 VDD vias_gen$15$1
X$28 VDD vias_gen$17$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1

.SUBCKT vias_gen$3 \$1
.ENDS vias_gen$3

.SUBCKT vias_gen$2 \$1
.ENDS vias_gen$2

.SUBCKT vias_gen \$1
.ENDS vias_gen

.SUBCKT rovcel2_LVT$2$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$25 OUT sky130_gnd nfet$3$2$1$1$1$1
X$2 GND GND \$28 OUT sky130_gnd nfet$3$2$1$1$1$1
X$3 IN OUT GND nfet$5$1$1$1$1
X$4 IN GND OUT nfet$5$1$1$1$1
X$5 GND vias_gen$17$2$1$1$1$1
X$6 GND vias_gen$17$2$1$1$1$1
X$7 GND vias_gen$15$2$1$1$1$1
X$8 OUT vias_gen$12$2$1$1$1$1
X$9 OUT vias_gen$8$2$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$2$1$1$1$1
X$11 VDD VDD \$28 OUT pfet$5$2$1$1$1$1
X$12 OUT vias_gen$8$2$1$1$1$1
X$13 OUT vias_gen$12$2$1$1$1$1
X$14 IN OUT VDD VDD pfet$4$2$1$1$1$1
X$15 IN VDD OUT VDD pfet$4$2$1$1$1$1
X$16 OUT vias_gen$13$2$1$1$1$1
X$17 IN VDD OUT VDD pfet$4$2$1$1$1$1
X$18 OUT vias_gen$13$2$1$1$1$1
X$19 IN OUT VDD VDD pfet$4$2$1$1$1$1
X$20 OUT vias_gen$16$2$1$1$1$1
X$21 OUT vias_gen$16$2$1$1$1$1
X$22 IN vias_gen$14$2$1$1$1$1
X$23 IN vias_gen$14$2$1$1$1$1
X$24 IN vias_gen$14$2$1$1$1$1
X$25 IN vias_gen$14$2$1$1$1$1
X$26 VDD vias_gen$17$2$1$1$1$1
X$27 VDD vias_gen$17$2$1$1$1$1
X$28 VDD vias_gen$15$2$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$2$1$1$1$1

.SUBCKT rovcel2_LVT$1$1$1$1$1$1 GND OUT IN VDD sky130_gnd
X$1 GND GND \$27 OUT sky130_gnd nfet$3$1$1$1$1$1$1
X$2 GND GND \$25 OUT sky130_gnd nfet$3$1$1$1$1$1$1
X$3 IN GND OUT nfet$4$1$1$1$1$1
X$4 GND vias_gen$17$1$1$1$1$1$1
X$5 GND vias_gen$15$1$1$1$1$1$1
X$6 GND vias_gen$17$1$1$1$1$1$1
X$7 IN OUT GND nfet$4$1$1$1$1$1
X$8 OUT vias_gen$12$1$1$1$1$1$1
X$9 OUT vias_gen$8$1$1$1$1$1$1
X$10 VDD VDD \$25 OUT pfet$5$1$1$1$1$1$1
X$11 VDD VDD \$27 OUT pfet$5$1$1$1$1$1$1
X$12 OUT vias_gen$8$1$1$1$1$1$1
X$13 OUT vias_gen$12$1$1$1$1$1$1
X$14 OUT vias_gen$16$1$1$1$1$1$1
X$15 OUT vias_gen$16$1$1$1$1$1$1
X$16 IN OUT VDD VDD pfet$4$1$1$1$1$1$1
X$17 OUT vias_gen$13$1$1$1$1$1$1
X$18 IN VDD OUT VDD pfet$4$1$1$1$1$1$1
X$19 OUT vias_gen$13$1$1$1$1$1$1
X$20 IN VDD OUT VDD pfet$4$1$1$1$1$1$1
X$21 IN OUT VDD VDD pfet$4$1$1$1$1$1$1
X$22 IN vias_gen$14$1$1$1$1$1$1
X$23 IN vias_gen$14$1$1$1$1$1$1
X$24 IN vias_gen$14$1$1$1$1$1$1
X$25 IN vias_gen$14$1$1$1$1$1$1
X$26 VDD vias_gen$17$1$1$1$1$1$1
X$27 VDD vias_gen$15$1$1$1$1$1$1
X$28 VDD vias_gen$17$1$1$1$1$1$1
M$1 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$3 VDD IN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=1.425 AD=0.7125
+ PS=10.1 PD=5.05
M$4 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 AS=0.7125 AD=1.425
+ PS=5.05 PD=10.1
M$5 OUT IN GND sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
M$6 GND IN OUT sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 AS=0.63
+ AD=0.63 PS=4.8 PD=4.8
.ENDS rovcel2_LVT$1$1$1$1$1$1

.SUBCKT vias_gen$8$2$1$1$1$1$1$1 \$1
.ENDS vias_gen$8$2$1$1$1$1$1$1

.SUBCKT vias_gen$13$2$1$1$1$1$1$1 \$1
.ENDS vias_gen$13$2$1$1$1$1$1$1

.SUBCKT vias_gen$12$2$1$1$1$1$1$1 \$1
.ENDS vias_gen$12$2$1$1$1$1$1$1

.SUBCKT vias_gen$14$2$1$1$1$1$1$1 \$1
.ENDS vias_gen$14$2$1$1$1$1$1$1

.SUBCKT pfet$4$2$1$1$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$1$1$1$1$1

.SUBCKT vias_gen$15$2$1$1$1$1$1$1 \$1
.ENDS vias_gen$15$2$1$1$1$1$1$1

.SUBCKT nfet$5$1$1$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$5$1$1$1$1$1$1

.SUBCKT vias_gen$16$2$1$1$1$1$1$1 \$1
.ENDS vias_gen$16$2$1$1$1$1$1$1

.SUBCKT vias_gen$17$2$1$1$1$1$1$1 \$1
.ENDS vias_gen$17$2$1$1$1$1$1$1

.SUBCKT pfet$5$2$1$1$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$1$1$1$1$1

.SUBCKT nfet$3$2$1$1$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$1$1$1$1$1

.SUBCKT nfet$3$1$1$1$1$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$16$1$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$16$1$1$1$1$1$1$1$1

.SUBCKT nfet$4$1$1$1$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$1$1$1$1$1$1

.SUBCKT vias_gen$15$1$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$15$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$14$1$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$14$1$1$1$1$1$1$1$1

.SUBCKT pfet$4$1$1$1$1$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$13$1$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$13$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$12$1$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$12$1$1$1$1$1$1$1$1

.SUBCKT pfet$5$1$1$1$1$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$8$1$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$8$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$17$1$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$17$1$1$1$1$1$1$1$1

.SUBCKT vias_gen$8$3$1$1$1$1$1 \$1
.ENDS vias_gen$8$3$1$1$1$1$1

.SUBCKT vias_gen$13$3$1$1$1$1$1 \$1
.ENDS vias_gen$13$3$1$1$1$1$1

.SUBCKT vias_gen$12$3$1$1$1$1$1 \$1
.ENDS vias_gen$12$3$1$1$1$1$1

.SUBCKT vias_gen$14$3$1$1$1$1$1 \$1
.ENDS vias_gen$14$3$1$1$1$1$1

.SUBCKT pfet$4$3$1$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$1$1$1$1$1

.SUBCKT vias_gen$15$3$1$1$1$1$1 \$1
.ENDS vias_gen$15$3$1$1$1$1$1

.SUBCKT nfet$6$1$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$6$1$1$1$1$1

.SUBCKT vias_gen$16$3$1$1$1$1$1 \$1
.ENDS vias_gen$16$3$1$1$1$1$1

.SUBCKT vias_gen$17$3$1$1$1$1$1 \$1
.ENDS vias_gen$17$3$1$1$1$1$1

.SUBCKT pfet$5$3$1$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$1$1$1$1$1

.SUBCKT nfet$3$3$1$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$1$1$1$1$1

.SUBCKT nfet$3$1$2$1$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$1$1$1$1$1

.SUBCKT vias_gen$16$1$2$1$1$1$1$1 \$1
.ENDS vias_gen$16$1$2$1$1$1$1$1

.SUBCKT nfet$4$2$1$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$2$1$1$1$1$1

.SUBCKT vias_gen$15$1$2$1$1$1$1$1 \$1
.ENDS vias_gen$15$1$2$1$1$1$1$1

.SUBCKT vias_gen$14$1$2$1$1$1$1$1 \$1
.ENDS vias_gen$14$1$2$1$1$1$1$1

.SUBCKT pfet$4$1$2$1$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$1$1$1$1$1

.SUBCKT vias_gen$13$1$2$1$1$1$1$1 \$1
.ENDS vias_gen$13$1$2$1$1$1$1$1

.SUBCKT vias_gen$12$1$2$1$1$1$1$1 \$1
.ENDS vias_gen$12$1$2$1$1$1$1$1

.SUBCKT pfet$5$1$2$1$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$1$1$1$1$1

.SUBCKT vias_gen$8$1$2$1$1$1$1$1 \$1
.ENDS vias_gen$8$1$2$1$1$1$1$1

.SUBCKT vias_gen$17$1$2$1$1$1$1$1 \$1
.ENDS vias_gen$17$1$2$1$1$1$1$1

.SUBCKT vias_gen$8$2$2$1$1$1$1 \$1
.ENDS vias_gen$8$2$2$1$1$1$1

.SUBCKT vias_gen$13$2$2$1$1$1$1 \$1
.ENDS vias_gen$13$2$2$1$1$1$1

.SUBCKT vias_gen$12$2$2$1$1$1$1 \$1
.ENDS vias_gen$12$2$2$1$1$1$1

.SUBCKT vias_gen$14$2$2$1$1$1$1 \$1
.ENDS vias_gen$14$2$2$1$1$1$1

.SUBCKT pfet$4$2$2$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$2$1$1$1$1

.SUBCKT vias_gen$15$2$2$1$1$1$1 \$1
.ENDS vias_gen$15$2$2$1$1$1$1

.SUBCKT nfet$5$2$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$5$2$1$1$1$1

.SUBCKT vias_gen$16$2$2$1$1$1$1 \$1
.ENDS vias_gen$16$2$2$1$1$1$1

.SUBCKT vias_gen$17$2$2$1$1$1$1 \$1
.ENDS vias_gen$17$2$2$1$1$1$1

.SUBCKT pfet$5$2$2$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$2$1$1$1$1

.SUBCKT nfet$3$2$2$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$2$1$1$1$1

.SUBCKT nfet$3$1$1$2$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$2$1$1$1$1

.SUBCKT vias_gen$16$1$1$2$1$1$1$1 \$1
.ENDS vias_gen$16$1$1$2$1$1$1$1

.SUBCKT nfet$4$1$2$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$2$1$1$1$1

.SUBCKT vias_gen$15$1$1$2$1$1$1$1 \$1
.ENDS vias_gen$15$1$1$2$1$1$1$1

.SUBCKT vias_gen$14$1$1$2$1$1$1$1 \$1
.ENDS vias_gen$14$1$1$2$1$1$1$1

.SUBCKT pfet$4$1$1$2$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$2$1$1$1$1

.SUBCKT vias_gen$13$1$1$2$1$1$1$1 \$1
.ENDS vias_gen$13$1$1$2$1$1$1$1

.SUBCKT vias_gen$12$1$1$2$1$1$1$1 \$1
.ENDS vias_gen$12$1$1$2$1$1$1$1

.SUBCKT pfet$5$1$1$2$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$2$1$1$1$1

.SUBCKT vias_gen$8$1$1$2$1$1$1$1 \$1
.ENDS vias_gen$8$1$1$2$1$1$1$1

.SUBCKT vias_gen$17$1$1$2$1$1$1$1 \$1
.ENDS vias_gen$17$1$1$2$1$1$1$1

.SUBCKT vias_gen$8$2$1$2$1$1$1 \$1
.ENDS vias_gen$8$2$1$2$1$1$1

.SUBCKT vias_gen$13$2$1$2$1$1$1 \$1
.ENDS vias_gen$13$2$1$2$1$1$1

.SUBCKT vias_gen$12$2$1$2$1$1$1 \$1
.ENDS vias_gen$12$2$1$2$1$1$1

.SUBCKT vias_gen$14$2$1$2$1$1$1 \$1
.ENDS vias_gen$14$2$1$2$1$1$1

.SUBCKT pfet$4$2$1$2$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$2$1$1$1

.SUBCKT vias_gen$15$2$1$2$1$1$1 \$1
.ENDS vias_gen$15$2$1$2$1$1$1

.SUBCKT nfet$5$1$2$1$1$1 \$1 \$2 \$3
.ENDS nfet$5$1$2$1$1$1

.SUBCKT vias_gen$16$2$1$2$1$1$1 \$1
.ENDS vias_gen$16$2$1$2$1$1$1

.SUBCKT vias_gen$17$2$1$2$1$1$1 \$1
.ENDS vias_gen$17$2$1$2$1$1$1

.SUBCKT pfet$5$2$1$2$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$2$1$1$1

.SUBCKT nfet$3$2$1$2$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$2$1$1$1

.SUBCKT nfet$3$1$1$1$2$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$2$1$1$1

.SUBCKT vias_gen$16$1$1$1$2$1$1$1 \$1
.ENDS vias_gen$16$1$1$1$2$1$1$1

.SUBCKT nfet$4$1$1$2$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$1$2$1$1$1

.SUBCKT vias_gen$15$1$1$1$2$1$1$1 \$1
.ENDS vias_gen$15$1$1$1$2$1$1$1

.SUBCKT vias_gen$14$1$1$1$2$1$1$1 \$1
.ENDS vias_gen$14$1$1$1$2$1$1$1

.SUBCKT pfet$4$1$1$1$2$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$2$1$1$1

.SUBCKT vias_gen$13$1$1$1$2$1$1$1 \$1
.ENDS vias_gen$13$1$1$1$2$1$1$1

.SUBCKT vias_gen$12$1$1$1$2$1$1$1 \$1
.ENDS vias_gen$12$1$1$1$2$1$1$1

.SUBCKT pfet$5$1$1$1$2$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$2$1$1$1

.SUBCKT vias_gen$8$1$1$1$2$1$1$1 \$1
.ENDS vias_gen$8$1$1$1$2$1$1$1

.SUBCKT vias_gen$17$1$1$1$2$1$1$1 \$1
.ENDS vias_gen$17$1$1$1$2$1$1$1

.SUBCKT vias_gen$8$3$2$1$1$1 \$1
.ENDS vias_gen$8$3$2$1$1$1

.SUBCKT vias_gen$13$3$2$1$1$1 \$1
.ENDS vias_gen$13$3$2$1$1$1

.SUBCKT vias_gen$12$3$2$1$1$1 \$1
.ENDS vias_gen$12$3$2$1$1$1

.SUBCKT vias_gen$14$3$2$1$1$1 \$1
.ENDS vias_gen$14$3$2$1$1$1

.SUBCKT pfet$4$3$2$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$2$1$1$1

.SUBCKT vias_gen$15$3$2$1$1$1 \$1
.ENDS vias_gen$15$3$2$1$1$1

.SUBCKT nfet$6$2$1$1$1 \$1 \$2 \$3
.ENDS nfet$6$2$1$1$1

.SUBCKT vias_gen$16$3$2$1$1$1 \$1
.ENDS vias_gen$16$3$2$1$1$1

.SUBCKT vias_gen$17$3$2$1$1$1 \$1
.ENDS vias_gen$17$3$2$1$1$1

.SUBCKT pfet$5$3$2$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$2$1$1$1

.SUBCKT nfet$3$3$2$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$2$1$1$1

.SUBCKT nfet$3$1$2$2$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$2$1$1$1

.SUBCKT vias_gen$16$1$2$2$1$1$1 \$1
.ENDS vias_gen$16$1$2$2$1$1$1

.SUBCKT nfet$4$2$2$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$2$2$1$1$1

.SUBCKT vias_gen$15$1$2$2$1$1$1 \$1
.ENDS vias_gen$15$1$2$2$1$1$1

.SUBCKT vias_gen$14$1$2$2$1$1$1 \$1
.ENDS vias_gen$14$1$2$2$1$1$1

.SUBCKT pfet$4$1$2$2$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$2$1$1$1

.SUBCKT vias_gen$13$1$2$2$1$1$1 \$1
.ENDS vias_gen$13$1$2$2$1$1$1

.SUBCKT vias_gen$12$1$2$2$1$1$1 \$1
.ENDS vias_gen$12$1$2$2$1$1$1

.SUBCKT pfet$5$1$2$2$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$2$1$1$1

.SUBCKT vias_gen$8$1$2$2$1$1$1 \$1
.ENDS vias_gen$8$1$2$2$1$1$1

.SUBCKT vias_gen$17$1$2$2$1$1$1 \$1
.ENDS vias_gen$17$1$2$2$1$1$1

.SUBCKT vias_gen$8$2$1$1$1$2$1 \$1
.ENDS vias_gen$8$2$1$1$1$2$1

.SUBCKT vias_gen$13$2$1$1$1$2$1 \$1
.ENDS vias_gen$13$2$1$1$1$2$1

.SUBCKT vias_gen$12$2$1$1$1$2$1 \$1
.ENDS vias_gen$12$2$1$1$1$2$1

.SUBCKT vias_gen$14$2$1$1$1$2$1 \$1
.ENDS vias_gen$14$2$1$1$1$2$1

.SUBCKT pfet$4$2$1$1$1$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$1$1$2$1

.SUBCKT vias_gen$15$2$1$1$1$2$1 \$1
.ENDS vias_gen$15$2$1$1$1$2$1

.SUBCKT nfet$5$1$1$1$2$1 \$1 \$2 \$3
.ENDS nfet$5$1$1$1$2$1

.SUBCKT vias_gen$16$2$1$1$1$2$1 \$1
.ENDS vias_gen$16$2$1$1$1$2$1

.SUBCKT vias_gen$17$2$1$1$1$2$1 \$1
.ENDS vias_gen$17$2$1$1$1$2$1

.SUBCKT pfet$5$2$1$1$1$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$1$1$2$1

.SUBCKT nfet$3$2$1$1$1$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$1$1$2$1

.SUBCKT nfet$3$1$1$1$1$1$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$1$1$2$1

.SUBCKT vias_gen$16$1$1$1$1$1$2$1 \$1
.ENDS vias_gen$16$1$1$1$1$1$2$1

.SUBCKT nfet$4$1$1$1$1$2$1 \$1 \$2 \$3
.ENDS nfet$4$1$1$1$1$2$1

.SUBCKT vias_gen$15$1$1$1$1$1$2$1 \$1
.ENDS vias_gen$15$1$1$1$1$1$2$1

.SUBCKT vias_gen$14$1$1$1$1$1$2$1 \$1
.ENDS vias_gen$14$1$1$1$1$1$2$1

.SUBCKT pfet$4$1$1$1$1$1$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$1$1$2$1

.SUBCKT vias_gen$13$1$1$1$1$1$2$1 \$1
.ENDS vias_gen$13$1$1$1$1$1$2$1

.SUBCKT vias_gen$12$1$1$1$1$1$2$1 \$1
.ENDS vias_gen$12$1$1$1$1$1$2$1

.SUBCKT pfet$5$1$1$1$1$1$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$1$1$2$1

.SUBCKT vias_gen$8$1$1$1$1$1$2$1 \$1
.ENDS vias_gen$8$1$1$1$1$1$2$1

.SUBCKT vias_gen$17$1$1$1$1$1$2$1 \$1
.ENDS vias_gen$17$1$1$1$1$1$2$1

.SUBCKT vias_gen$8$3$1$1$2$1 \$1
.ENDS vias_gen$8$3$1$1$2$1

.SUBCKT vias_gen$13$3$1$1$2$1 \$1
.ENDS vias_gen$13$3$1$1$2$1

.SUBCKT vias_gen$12$3$1$1$2$1 \$1
.ENDS vias_gen$12$3$1$1$2$1

.SUBCKT vias_gen$14$3$1$1$2$1 \$1
.ENDS vias_gen$14$3$1$1$2$1

.SUBCKT pfet$4$3$1$1$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$1$1$2$1

.SUBCKT vias_gen$15$3$1$1$2$1 \$1
.ENDS vias_gen$15$3$1$1$2$1

.SUBCKT nfet$6$1$1$2$1 \$1 \$2 \$3
.ENDS nfet$6$1$1$2$1

.SUBCKT vias_gen$16$3$1$1$2$1 \$1
.ENDS vias_gen$16$3$1$1$2$1

.SUBCKT vias_gen$17$3$1$1$2$1 \$1
.ENDS vias_gen$17$3$1$1$2$1

.SUBCKT pfet$5$3$1$1$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$1$1$2$1

.SUBCKT nfet$3$3$1$1$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$1$1$2$1

.SUBCKT nfet$3$1$2$1$1$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$1$1$2$1

.SUBCKT vias_gen$16$1$2$1$1$2$1 \$1
.ENDS vias_gen$16$1$2$1$1$2$1

.SUBCKT nfet$4$2$1$1$2$1 \$1 \$2 \$3
.ENDS nfet$4$2$1$1$2$1

.SUBCKT vias_gen$15$1$2$1$1$2$1 \$1
.ENDS vias_gen$15$1$2$1$1$2$1

.SUBCKT vias_gen$14$1$2$1$1$2$1 \$1
.ENDS vias_gen$14$1$2$1$1$2$1

.SUBCKT pfet$4$1$2$1$1$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$1$1$2$1

.SUBCKT vias_gen$13$1$2$1$1$2$1 \$1
.ENDS vias_gen$13$1$2$1$1$2$1

.SUBCKT vias_gen$12$1$2$1$1$2$1 \$1
.ENDS vias_gen$12$1$2$1$1$2$1

.SUBCKT pfet$5$1$2$1$1$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$1$1$2$1

.SUBCKT vias_gen$8$1$2$1$1$2$1 \$1
.ENDS vias_gen$8$1$2$1$1$2$1

.SUBCKT vias_gen$17$1$2$1$1$2$1 \$1
.ENDS vias_gen$17$1$2$1$1$2$1

.SUBCKT vias_gen$8$2$2$1$2$1 \$1
.ENDS vias_gen$8$2$2$1$2$1

.SUBCKT vias_gen$13$2$2$1$2$1 \$1
.ENDS vias_gen$13$2$2$1$2$1

.SUBCKT vias_gen$12$2$2$1$2$1 \$1
.ENDS vias_gen$12$2$2$1$2$1

.SUBCKT vias_gen$14$2$2$1$2$1 \$1
.ENDS vias_gen$14$2$2$1$2$1

.SUBCKT pfet$4$2$2$1$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$2$1$2$1

.SUBCKT vias_gen$15$2$2$1$2$1 \$1
.ENDS vias_gen$15$2$2$1$2$1

.SUBCKT nfet$5$2$1$2$1 \$1 \$2 \$3
.ENDS nfet$5$2$1$2$1

.SUBCKT vias_gen$16$2$2$1$2$1 \$1
.ENDS vias_gen$16$2$2$1$2$1

.SUBCKT vias_gen$17$2$2$1$2$1 \$1
.ENDS vias_gen$17$2$2$1$2$1

.SUBCKT pfet$5$2$2$1$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$2$1$2$1

.SUBCKT nfet$3$2$2$1$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$2$1$2$1

.SUBCKT nfet$3$1$1$2$1$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$2$1$2$1

.SUBCKT vias_gen$16$1$1$2$1$2$1 \$1
.ENDS vias_gen$16$1$1$2$1$2$1

.SUBCKT nfet$4$1$2$1$2$1 \$1 \$2 \$3
.ENDS nfet$4$1$2$1$2$1

.SUBCKT vias_gen$15$1$1$2$1$2$1 \$1
.ENDS vias_gen$15$1$1$2$1$2$1

.SUBCKT vias_gen$14$1$1$2$1$2$1 \$1
.ENDS vias_gen$14$1$1$2$1$2$1

.SUBCKT pfet$4$1$1$2$1$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$2$1$2$1

.SUBCKT vias_gen$13$1$1$2$1$2$1 \$1
.ENDS vias_gen$13$1$1$2$1$2$1

.SUBCKT vias_gen$12$1$1$2$1$2$1 \$1
.ENDS vias_gen$12$1$1$2$1$2$1

.SUBCKT pfet$5$1$1$2$1$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$2$1$2$1

.SUBCKT vias_gen$8$1$1$2$1$2$1 \$1
.ENDS vias_gen$8$1$1$2$1$2$1

.SUBCKT vias_gen$17$1$1$2$1$2$1 \$1
.ENDS vias_gen$17$1$1$2$1$2$1

.SUBCKT vias_gen$8$2$1$2$2$1 \$1
.ENDS vias_gen$8$2$1$2$2$1

.SUBCKT vias_gen$13$2$1$2$2$1 \$1
.ENDS vias_gen$13$2$1$2$2$1

.SUBCKT vias_gen$12$2$1$2$2$1 \$1
.ENDS vias_gen$12$2$1$2$2$1

.SUBCKT vias_gen$14$2$1$2$2$1 \$1
.ENDS vias_gen$14$2$1$2$2$1

.SUBCKT pfet$4$2$1$2$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$2$2$1

.SUBCKT vias_gen$15$2$1$2$2$1 \$1
.ENDS vias_gen$15$2$1$2$2$1

.SUBCKT nfet$5$1$2$2$1 \$1 \$2 \$3
.ENDS nfet$5$1$2$2$1

.SUBCKT vias_gen$16$2$1$2$2$1 \$1
.ENDS vias_gen$16$2$1$2$2$1

.SUBCKT vias_gen$17$2$1$2$2$1 \$1
.ENDS vias_gen$17$2$1$2$2$1

.SUBCKT pfet$5$2$1$2$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$2$2$1

.SUBCKT nfet$3$2$1$2$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$2$2$1

.SUBCKT nfet$3$1$1$1$2$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$2$2$1

.SUBCKT vias_gen$16$1$1$1$2$2$1 \$1
.ENDS vias_gen$16$1$1$1$2$2$1

.SUBCKT nfet$4$1$1$2$2$1 \$1 \$2 \$3
.ENDS nfet$4$1$1$2$2$1

.SUBCKT vias_gen$15$1$1$1$2$2$1 \$1
.ENDS vias_gen$15$1$1$1$2$2$1

.SUBCKT vias_gen$14$1$1$1$2$2$1 \$1
.ENDS vias_gen$14$1$1$1$2$2$1

.SUBCKT pfet$4$1$1$1$2$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$2$2$1

.SUBCKT vias_gen$13$1$1$1$2$2$1 \$1
.ENDS vias_gen$13$1$1$1$2$2$1

.SUBCKT vias_gen$12$1$1$1$2$2$1 \$1
.ENDS vias_gen$12$1$1$1$2$2$1

.SUBCKT pfet$5$1$1$1$2$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$2$2$1

.SUBCKT vias_gen$8$1$1$1$2$2$1 \$1
.ENDS vias_gen$8$1$1$1$2$2$1

.SUBCKT vias_gen$17$1$1$1$2$2$1 \$1
.ENDS vias_gen$17$1$1$1$2$2$1

.SUBCKT vias_gen$8$3$2$2$1 \$1
.ENDS vias_gen$8$3$2$2$1

.SUBCKT vias_gen$13$3$2$2$1 \$1
.ENDS vias_gen$13$3$2$2$1

.SUBCKT vias_gen$12$3$2$2$1 \$1
.ENDS vias_gen$12$3$2$2$1

.SUBCKT vias_gen$14$3$2$2$1 \$1
.ENDS vias_gen$14$3$2$2$1

.SUBCKT pfet$4$3$2$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$2$2$1

.SUBCKT vias_gen$15$3$2$2$1 \$1
.ENDS vias_gen$15$3$2$2$1

.SUBCKT nfet$6$2$2$1 \$1 \$2 \$3
.ENDS nfet$6$2$2$1

.SUBCKT vias_gen$16$3$2$2$1 \$1
.ENDS vias_gen$16$3$2$2$1

.SUBCKT vias_gen$17$3$2$2$1 \$1
.ENDS vias_gen$17$3$2$2$1

.SUBCKT pfet$5$3$2$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$2$2$1

.SUBCKT nfet$3$3$2$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$2$2$1

.SUBCKT nfet$3$1$2$2$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$2$2$1

.SUBCKT vias_gen$16$1$2$2$2$1 \$1
.ENDS vias_gen$16$1$2$2$2$1

.SUBCKT nfet$4$2$2$2$1 \$1 \$2 \$3
.ENDS nfet$4$2$2$2$1

.SUBCKT vias_gen$15$1$2$2$2$1 \$1
.ENDS vias_gen$15$1$2$2$2$1

.SUBCKT vias_gen$14$1$2$2$2$1 \$1
.ENDS vias_gen$14$1$2$2$2$1

.SUBCKT pfet$4$1$2$2$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$2$2$1

.SUBCKT vias_gen$13$1$2$2$2$1 \$1
.ENDS vias_gen$13$1$2$2$2$1

.SUBCKT vias_gen$12$1$2$2$2$1 \$1
.ENDS vias_gen$12$1$2$2$2$1

.SUBCKT pfet$5$1$2$2$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$2$2$1

.SUBCKT vias_gen$8$1$2$2$2$1 \$1
.ENDS vias_gen$8$1$2$2$2$1

.SUBCKT vias_gen$17$1$2$2$2$1 \$1
.ENDS vias_gen$17$1$2$2$2$1

.SUBCKT vias_gen$8$2$1$1$1$1$2 \$1
.ENDS vias_gen$8$2$1$1$1$1$2

.SUBCKT vias_gen$13$2$1$1$1$1$2 \$1
.ENDS vias_gen$13$2$1$1$1$1$2

.SUBCKT vias_gen$12$2$1$1$1$1$2 \$1
.ENDS vias_gen$12$2$1$1$1$1$2

.SUBCKT vias_gen$14$2$1$1$1$1$2 \$1
.ENDS vias_gen$14$2$1$1$1$1$2

.SUBCKT pfet$4$2$1$1$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$1$1$1$2

.SUBCKT vias_gen$15$2$1$1$1$1$2 \$1
.ENDS vias_gen$15$2$1$1$1$1$2

.SUBCKT nfet$5$1$1$1$1$2 \$1 \$2 \$3
.ENDS nfet$5$1$1$1$1$2

.SUBCKT vias_gen$16$2$1$1$1$1$2 \$1
.ENDS vias_gen$16$2$1$1$1$1$2

.SUBCKT vias_gen$17$2$1$1$1$1$2 \$1
.ENDS vias_gen$17$2$1$1$1$1$2

.SUBCKT pfet$5$2$1$1$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$1$1$1$2

.SUBCKT nfet$3$2$1$1$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$1$1$1$2

.SUBCKT nfet$3$1$1$1$1$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$1$1$1$2

.SUBCKT vias_gen$16$1$1$1$1$1$1$2 \$1
.ENDS vias_gen$16$1$1$1$1$1$1$2

.SUBCKT nfet$4$1$1$1$1$1$2 \$1 \$2 \$3
.ENDS nfet$4$1$1$1$1$1$2

.SUBCKT vias_gen$15$1$1$1$1$1$1$2 \$1
.ENDS vias_gen$15$1$1$1$1$1$1$2

.SUBCKT vias_gen$14$1$1$1$1$1$1$2 \$1
.ENDS vias_gen$14$1$1$1$1$1$1$2

.SUBCKT pfet$4$1$1$1$1$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$1$1$1$2

.SUBCKT vias_gen$13$1$1$1$1$1$1$2 \$1
.ENDS vias_gen$13$1$1$1$1$1$1$2

.SUBCKT vias_gen$12$1$1$1$1$1$1$2 \$1
.ENDS vias_gen$12$1$1$1$1$1$1$2

.SUBCKT pfet$5$1$1$1$1$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$1$1$1$2

.SUBCKT vias_gen$8$1$1$1$1$1$1$2 \$1
.ENDS vias_gen$8$1$1$1$1$1$1$2

.SUBCKT vias_gen$17$1$1$1$1$1$1$2 \$1
.ENDS vias_gen$17$1$1$1$1$1$1$2

.SUBCKT vias_gen$8$3$1$1$1$2 \$1
.ENDS vias_gen$8$3$1$1$1$2

.SUBCKT vias_gen$13$3$1$1$1$2 \$1
.ENDS vias_gen$13$3$1$1$1$2

.SUBCKT vias_gen$12$3$1$1$1$2 \$1
.ENDS vias_gen$12$3$1$1$1$2

.SUBCKT vias_gen$14$3$1$1$1$2 \$1
.ENDS vias_gen$14$3$1$1$1$2

.SUBCKT pfet$4$3$1$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$1$1$1$2

.SUBCKT vias_gen$15$3$1$1$1$2 \$1
.ENDS vias_gen$15$3$1$1$1$2

.SUBCKT nfet$6$1$1$1$2 \$1 \$2 \$3
.ENDS nfet$6$1$1$1$2

.SUBCKT vias_gen$16$3$1$1$1$2 \$1
.ENDS vias_gen$16$3$1$1$1$2

.SUBCKT vias_gen$17$3$1$1$1$2 \$1
.ENDS vias_gen$17$3$1$1$1$2

.SUBCKT pfet$5$3$1$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$1$1$1$2

.SUBCKT nfet$3$3$1$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$1$1$1$2

.SUBCKT nfet$3$1$2$1$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$1$1$1$2

.SUBCKT vias_gen$16$1$2$1$1$1$2 \$1
.ENDS vias_gen$16$1$2$1$1$1$2

.SUBCKT nfet$4$2$1$1$1$2 \$1 \$2 \$3
.ENDS nfet$4$2$1$1$1$2

.SUBCKT vias_gen$15$1$2$1$1$1$2 \$1
.ENDS vias_gen$15$1$2$1$1$1$2

.SUBCKT vias_gen$14$1$2$1$1$1$2 \$1
.ENDS vias_gen$14$1$2$1$1$1$2

.SUBCKT pfet$4$1$2$1$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$1$1$1$2

.SUBCKT vias_gen$13$1$2$1$1$1$2 \$1
.ENDS vias_gen$13$1$2$1$1$1$2

.SUBCKT vias_gen$12$1$2$1$1$1$2 \$1
.ENDS vias_gen$12$1$2$1$1$1$2

.SUBCKT pfet$5$1$2$1$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$1$1$1$2

.SUBCKT vias_gen$8$1$2$1$1$1$2 \$1
.ENDS vias_gen$8$1$2$1$1$1$2

.SUBCKT vias_gen$17$1$2$1$1$1$2 \$1
.ENDS vias_gen$17$1$2$1$1$1$2

.SUBCKT vias_gen$8$2$2$1$1$2 \$1
.ENDS vias_gen$8$2$2$1$1$2

.SUBCKT vias_gen$13$2$2$1$1$2 \$1
.ENDS vias_gen$13$2$2$1$1$2

.SUBCKT vias_gen$12$2$2$1$1$2 \$1
.ENDS vias_gen$12$2$2$1$1$2

.SUBCKT vias_gen$14$2$2$1$1$2 \$1
.ENDS vias_gen$14$2$2$1$1$2

.SUBCKT pfet$4$2$2$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$2$1$1$2

.SUBCKT vias_gen$15$2$2$1$1$2 \$1
.ENDS vias_gen$15$2$2$1$1$2

.SUBCKT nfet$5$2$1$1$2 \$1 \$2 \$3
.ENDS nfet$5$2$1$1$2

.SUBCKT vias_gen$16$2$2$1$1$2 \$1
.ENDS vias_gen$16$2$2$1$1$2

.SUBCKT vias_gen$17$2$2$1$1$2 \$1
.ENDS vias_gen$17$2$2$1$1$2

.SUBCKT pfet$5$2$2$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$2$1$1$2

.SUBCKT nfet$3$2$2$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$2$1$1$2

.SUBCKT nfet$3$1$1$2$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$2$1$1$2

.SUBCKT vias_gen$16$1$1$2$1$1$2 \$1
.ENDS vias_gen$16$1$1$2$1$1$2

.SUBCKT nfet$4$1$2$1$1$2 \$1 \$2 \$3
.ENDS nfet$4$1$2$1$1$2

.SUBCKT vias_gen$15$1$1$2$1$1$2 \$1
.ENDS vias_gen$15$1$1$2$1$1$2

.SUBCKT vias_gen$14$1$1$2$1$1$2 \$1
.ENDS vias_gen$14$1$1$2$1$1$2

.SUBCKT pfet$4$1$1$2$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$2$1$1$2

.SUBCKT vias_gen$13$1$1$2$1$1$2 \$1
.ENDS vias_gen$13$1$1$2$1$1$2

.SUBCKT vias_gen$12$1$1$2$1$1$2 \$1
.ENDS vias_gen$12$1$1$2$1$1$2

.SUBCKT pfet$5$1$1$2$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$2$1$1$2

.SUBCKT vias_gen$8$1$1$2$1$1$2 \$1
.ENDS vias_gen$8$1$1$2$1$1$2

.SUBCKT vias_gen$17$1$1$2$1$1$2 \$1
.ENDS vias_gen$17$1$1$2$1$1$2

.SUBCKT vias_gen$8$2$1$2$1$2 \$1
.ENDS vias_gen$8$2$1$2$1$2

.SUBCKT vias_gen$13$2$1$2$1$2 \$1
.ENDS vias_gen$13$2$1$2$1$2

.SUBCKT vias_gen$12$2$1$2$1$2 \$1
.ENDS vias_gen$12$2$1$2$1$2

.SUBCKT vias_gen$14$2$1$2$1$2 \$1
.ENDS vias_gen$14$2$1$2$1$2

.SUBCKT pfet$4$2$1$2$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$2$1$2

.SUBCKT vias_gen$15$2$1$2$1$2 \$1
.ENDS vias_gen$15$2$1$2$1$2

.SUBCKT nfet$5$1$2$1$2 \$1 \$2 \$3
.ENDS nfet$5$1$2$1$2

.SUBCKT vias_gen$16$2$1$2$1$2 \$1
.ENDS vias_gen$16$2$1$2$1$2

.SUBCKT vias_gen$17$2$1$2$1$2 \$1
.ENDS vias_gen$17$2$1$2$1$2

.SUBCKT pfet$5$2$1$2$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$2$1$2

.SUBCKT nfet$3$2$1$2$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$2$1$2

.SUBCKT nfet$3$1$1$1$2$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$2$1$2

.SUBCKT vias_gen$16$1$1$1$2$1$2 \$1
.ENDS vias_gen$16$1$1$1$2$1$2

.SUBCKT nfet$4$1$1$2$1$2 \$1 \$2 \$3
.ENDS nfet$4$1$1$2$1$2

.SUBCKT vias_gen$15$1$1$1$2$1$2 \$1
.ENDS vias_gen$15$1$1$1$2$1$2

.SUBCKT vias_gen$14$1$1$1$2$1$2 \$1
.ENDS vias_gen$14$1$1$1$2$1$2

.SUBCKT pfet$4$1$1$1$2$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$2$1$2

.SUBCKT vias_gen$13$1$1$1$2$1$2 \$1
.ENDS vias_gen$13$1$1$1$2$1$2

.SUBCKT vias_gen$12$1$1$1$2$1$2 \$1
.ENDS vias_gen$12$1$1$1$2$1$2

.SUBCKT pfet$5$1$1$1$2$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$2$1$2

.SUBCKT vias_gen$8$1$1$1$2$1$2 \$1
.ENDS vias_gen$8$1$1$1$2$1$2

.SUBCKT vias_gen$17$1$1$1$2$1$2 \$1
.ENDS vias_gen$17$1$1$1$2$1$2

.SUBCKT vias_gen$8$3$2$1$2 \$1
.ENDS vias_gen$8$3$2$1$2

.SUBCKT vias_gen$13$3$2$1$2 \$1
.ENDS vias_gen$13$3$2$1$2

.SUBCKT vias_gen$12$3$2$1$2 \$1
.ENDS vias_gen$12$3$2$1$2

.SUBCKT vias_gen$14$3$2$1$2 \$1
.ENDS vias_gen$14$3$2$1$2

.SUBCKT pfet$4$3$2$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$2$1$2

.SUBCKT vias_gen$15$3$2$1$2 \$1
.ENDS vias_gen$15$3$2$1$2

.SUBCKT nfet$6$2$1$2 \$1 \$2 \$3
.ENDS nfet$6$2$1$2

.SUBCKT vias_gen$16$3$2$1$2 \$1
.ENDS vias_gen$16$3$2$1$2

.SUBCKT vias_gen$17$3$2$1$2 \$1
.ENDS vias_gen$17$3$2$1$2

.SUBCKT pfet$5$3$2$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$2$1$2

.SUBCKT nfet$3$3$2$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$2$1$2

.SUBCKT nfet$3$1$2$2$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$2$1$2

.SUBCKT vias_gen$16$1$2$2$1$2 \$1
.ENDS vias_gen$16$1$2$2$1$2

.SUBCKT nfet$4$2$2$1$2 \$1 \$2 \$3
.ENDS nfet$4$2$2$1$2

.SUBCKT vias_gen$15$1$2$2$1$2 \$1
.ENDS vias_gen$15$1$2$2$1$2

.SUBCKT vias_gen$14$1$2$2$1$2 \$1
.ENDS vias_gen$14$1$2$2$1$2

.SUBCKT pfet$4$1$2$2$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$2$1$2

.SUBCKT vias_gen$13$1$2$2$1$2 \$1
.ENDS vias_gen$13$1$2$2$1$2

.SUBCKT vias_gen$12$1$2$2$1$2 \$1
.ENDS vias_gen$12$1$2$2$1$2

.SUBCKT pfet$5$1$2$2$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$2$1$2

.SUBCKT vias_gen$8$1$2$2$1$2 \$1
.ENDS vias_gen$8$1$2$2$1$2

.SUBCKT vias_gen$17$1$2$2$1$2 \$1
.ENDS vias_gen$17$1$2$2$1$2

.SUBCKT vias_gen$8$2$1$1$1$3 \$1
.ENDS vias_gen$8$2$1$1$1$3

.SUBCKT vias_gen$13$2$1$1$1$3 \$1
.ENDS vias_gen$13$2$1$1$1$3

.SUBCKT vias_gen$12$2$1$1$1$3 \$1
.ENDS vias_gen$12$2$1$1$1$3

.SUBCKT vias_gen$14$2$1$1$1$3 \$1
.ENDS vias_gen$14$2$1$1$1$3

.SUBCKT pfet$4$2$1$1$1$3 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$1$1$3

.SUBCKT vias_gen$15$2$1$1$1$3 \$1
.ENDS vias_gen$15$2$1$1$1$3

.SUBCKT nfet$5$1$1$1$3 \$1 \$2 \$3
.ENDS nfet$5$1$1$1$3

.SUBCKT vias_gen$16$2$1$1$1$3 \$1
.ENDS vias_gen$16$2$1$1$1$3

.SUBCKT vias_gen$17$2$1$1$1$3 \$1
.ENDS vias_gen$17$2$1$1$1$3

.SUBCKT pfet$5$2$1$1$1$3 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$1$1$3

.SUBCKT nfet$3$2$1$1$1$3 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$1$1$3

.SUBCKT nfet$3$1$1$1$1$1$3 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$1$1$3

.SUBCKT vias_gen$16$1$1$1$1$1$3 \$1
.ENDS vias_gen$16$1$1$1$1$1$3

.SUBCKT nfet$4$1$1$1$1$3 \$1 \$2 \$3
.ENDS nfet$4$1$1$1$1$3

.SUBCKT vias_gen$15$1$1$1$1$1$3 \$1
.ENDS vias_gen$15$1$1$1$1$1$3

.SUBCKT vias_gen$14$1$1$1$1$1$3 \$1
.ENDS vias_gen$14$1$1$1$1$1$3

.SUBCKT pfet$4$1$1$1$1$1$3 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$1$1$3

.SUBCKT vias_gen$13$1$1$1$1$1$3 \$1
.ENDS vias_gen$13$1$1$1$1$1$3

.SUBCKT vias_gen$12$1$1$1$1$1$3 \$1
.ENDS vias_gen$12$1$1$1$1$1$3

.SUBCKT pfet$5$1$1$1$1$1$3 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$1$1$3

.SUBCKT vias_gen$8$1$1$1$1$1$3 \$1
.ENDS vias_gen$8$1$1$1$1$1$3

.SUBCKT vias_gen$17$1$1$1$1$1$3 \$1
.ENDS vias_gen$17$1$1$1$1$1$3

.SUBCKT vias_gen$8$3$1$1$3 \$1
.ENDS vias_gen$8$3$1$1$3

.SUBCKT vias_gen$13$3$1$1$3 \$1
.ENDS vias_gen$13$3$1$1$3

.SUBCKT vias_gen$12$3$1$1$3 \$1
.ENDS vias_gen$12$3$1$1$3

.SUBCKT vias_gen$14$3$1$1$3 \$1
.ENDS vias_gen$14$3$1$1$3

.SUBCKT pfet$4$3$1$1$3 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$1$1$3

.SUBCKT vias_gen$15$3$1$1$3 \$1
.ENDS vias_gen$15$3$1$1$3

.SUBCKT nfet$6$1$1$3 \$1 \$2 \$3
.ENDS nfet$6$1$1$3

.SUBCKT vias_gen$16$3$1$1$3 \$1
.ENDS vias_gen$16$3$1$1$3

.SUBCKT vias_gen$17$3$1$1$3 \$1
.ENDS vias_gen$17$3$1$1$3

.SUBCKT pfet$5$3$1$1$3 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$1$1$3

.SUBCKT nfet$3$3$1$1$3 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$1$1$3

.SUBCKT nfet$3$1$2$1$1$3 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$1$1$3

.SUBCKT vias_gen$16$1$2$1$1$3 \$1
.ENDS vias_gen$16$1$2$1$1$3

.SUBCKT nfet$4$2$1$1$3 \$1 \$2 \$3
.ENDS nfet$4$2$1$1$3

.SUBCKT vias_gen$15$1$2$1$1$3 \$1
.ENDS vias_gen$15$1$2$1$1$3

.SUBCKT vias_gen$14$1$2$1$1$3 \$1
.ENDS vias_gen$14$1$2$1$1$3

.SUBCKT pfet$4$1$2$1$1$3 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$1$1$3

.SUBCKT vias_gen$13$1$2$1$1$3 \$1
.ENDS vias_gen$13$1$2$1$1$3

.SUBCKT vias_gen$12$1$2$1$1$3 \$1
.ENDS vias_gen$12$1$2$1$1$3

.SUBCKT pfet$5$1$2$1$1$3 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$1$1$3

.SUBCKT vias_gen$8$1$2$1$1$3 \$1
.ENDS vias_gen$8$1$2$1$1$3

.SUBCKT vias_gen$17$1$2$1$1$3 \$1
.ENDS vias_gen$17$1$2$1$1$3

.SUBCKT vias_gen$8$2$1$1$1$1$1 \$1
.ENDS vias_gen$8$2$1$1$1$1$1

.SUBCKT vias_gen$13$2$1$1$1$1$1 \$1
.ENDS vias_gen$13$2$1$1$1$1$1

.SUBCKT vias_gen$12$2$1$1$1$1$1 \$1
.ENDS vias_gen$12$2$1$1$1$1$1

.SUBCKT vias_gen$14$2$1$1$1$1$1 \$1
.ENDS vias_gen$14$2$1$1$1$1$1

.SUBCKT pfet$4$2$1$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$1$1$1$1

.SUBCKT vias_gen$15$2$1$1$1$1$1 \$1
.ENDS vias_gen$15$2$1$1$1$1$1

.SUBCKT nfet$5$1$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$5$1$1$1$1$1

.SUBCKT vias_gen$16$2$1$1$1$1$1 \$1
.ENDS vias_gen$16$2$1$1$1$1$1

.SUBCKT vias_gen$17$2$1$1$1$1$1 \$1
.ENDS vias_gen$17$2$1$1$1$1$1

.SUBCKT pfet$5$2$1$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$1$1$1$1

.SUBCKT nfet$3$2$1$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$1$1$1$1

.SUBCKT nfet$3$1$1$1$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$1$1$1$1

.SUBCKT vias_gen$16$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$16$1$1$1$1$1$1$1

.SUBCKT nfet$4$1$1$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$1$1$1$1$1

.SUBCKT vias_gen$15$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$15$1$1$1$1$1$1$1

.SUBCKT vias_gen$14$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$14$1$1$1$1$1$1$1

.SUBCKT pfet$4$1$1$1$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$1$1$1$1

.SUBCKT vias_gen$13$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$13$1$1$1$1$1$1$1

.SUBCKT vias_gen$12$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$12$1$1$1$1$1$1$1

.SUBCKT pfet$5$1$1$1$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$1$1$1$1

.SUBCKT vias_gen$8$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$8$1$1$1$1$1$1$1

.SUBCKT vias_gen$17$1$1$1$1$1$1$1 \$1
.ENDS vias_gen$17$1$1$1$1$1$1$1

.SUBCKT vias_gen$8$3$1$1$1$1 \$1
.ENDS vias_gen$8$3$1$1$1$1

.SUBCKT vias_gen$13$3$1$1$1$1 \$1
.ENDS vias_gen$13$3$1$1$1$1

.SUBCKT vias_gen$12$3$1$1$1$1 \$1
.ENDS vias_gen$12$3$1$1$1$1

.SUBCKT vias_gen$14$3$1$1$1$1 \$1
.ENDS vias_gen$14$3$1$1$1$1

.SUBCKT pfet$4$3$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$1$1$1$1

.SUBCKT vias_gen$15$3$1$1$1$1 \$1
.ENDS vias_gen$15$3$1$1$1$1

.SUBCKT nfet$6$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$6$1$1$1$1

.SUBCKT vias_gen$16$3$1$1$1$1 \$1
.ENDS vias_gen$16$3$1$1$1$1

.SUBCKT vias_gen$17$3$1$1$1$1 \$1
.ENDS vias_gen$17$3$1$1$1$1

.SUBCKT pfet$5$3$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$1$1$1$1

.SUBCKT nfet$3$3$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$1$1$1$1

.SUBCKT nfet$3$1$2$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$1$1$1$1

.SUBCKT vias_gen$16$1$2$1$1$1$1 \$1
.ENDS vias_gen$16$1$2$1$1$1$1

.SUBCKT nfet$4$2$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$2$1$1$1$1

.SUBCKT vias_gen$15$1$2$1$1$1$1 \$1
.ENDS vias_gen$15$1$2$1$1$1$1

.SUBCKT vias_gen$14$1$2$1$1$1$1 \$1
.ENDS vias_gen$14$1$2$1$1$1$1

.SUBCKT pfet$4$1$2$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$1$1$1$1

.SUBCKT vias_gen$13$1$2$1$1$1$1 \$1
.ENDS vias_gen$13$1$2$1$1$1$1

.SUBCKT vias_gen$12$1$2$1$1$1$1 \$1
.ENDS vias_gen$12$1$2$1$1$1$1

.SUBCKT pfet$5$1$2$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$1$1$1$1

.SUBCKT vias_gen$8$1$2$1$1$1$1 \$1
.ENDS vias_gen$8$1$2$1$1$1$1

.SUBCKT vias_gen$17$1$2$1$1$1$1 \$1
.ENDS vias_gen$17$1$2$1$1$1$1

.SUBCKT vias_gen$8$2$2$1$1$1 \$1
.ENDS vias_gen$8$2$2$1$1$1

.SUBCKT vias_gen$13$2$2$1$1$1 \$1
.ENDS vias_gen$13$2$2$1$1$1

.SUBCKT vias_gen$12$2$2$1$1$1 \$1
.ENDS vias_gen$12$2$2$1$1$1

.SUBCKT vias_gen$14$2$2$1$1$1 \$1
.ENDS vias_gen$14$2$2$1$1$1

.SUBCKT pfet$4$2$2$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$2$1$1$1

.SUBCKT vias_gen$15$2$2$1$1$1 \$1
.ENDS vias_gen$15$2$2$1$1$1

.SUBCKT nfet$5$2$1$1$1 \$1 \$2 \$3
.ENDS nfet$5$2$1$1$1

.SUBCKT vias_gen$16$2$2$1$1$1 \$1
.ENDS vias_gen$16$2$2$1$1$1

.SUBCKT vias_gen$17$2$2$1$1$1 \$1
.ENDS vias_gen$17$2$2$1$1$1

.SUBCKT pfet$5$2$2$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$2$1$1$1

.SUBCKT nfet$3$2$2$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$2$1$1$1

.SUBCKT nfet$3$1$1$2$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$2$1$1$1

.SUBCKT vias_gen$16$1$1$2$1$1$1 \$1
.ENDS vias_gen$16$1$1$2$1$1$1

.SUBCKT nfet$4$1$2$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$2$1$1$1

.SUBCKT vias_gen$15$1$1$2$1$1$1 \$1
.ENDS vias_gen$15$1$1$2$1$1$1

.SUBCKT vias_gen$14$1$1$2$1$1$1 \$1
.ENDS vias_gen$14$1$1$2$1$1$1

.SUBCKT pfet$4$1$1$2$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$2$1$1$1

.SUBCKT vias_gen$13$1$1$2$1$1$1 \$1
.ENDS vias_gen$13$1$1$2$1$1$1

.SUBCKT vias_gen$12$1$1$2$1$1$1 \$1
.ENDS vias_gen$12$1$1$2$1$1$1

.SUBCKT pfet$5$1$1$2$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$2$1$1$1

.SUBCKT vias_gen$8$1$1$2$1$1$1 \$1
.ENDS vias_gen$8$1$1$2$1$1$1

.SUBCKT vias_gen$17$1$1$2$1$1$1 \$1
.ENDS vias_gen$17$1$1$2$1$1$1

.SUBCKT vias_gen$8$2$1$2$1$1 \$1
.ENDS vias_gen$8$2$1$2$1$1

.SUBCKT vias_gen$13$2$1$2$1$1 \$1
.ENDS vias_gen$13$2$1$2$1$1

.SUBCKT vias_gen$12$2$1$2$1$1 \$1
.ENDS vias_gen$12$2$1$2$1$1

.SUBCKT vias_gen$14$2$1$2$1$1 \$1
.ENDS vias_gen$14$2$1$2$1$1

.SUBCKT pfet$4$2$1$2$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$2$1$1

.SUBCKT vias_gen$15$2$1$2$1$1 \$1
.ENDS vias_gen$15$2$1$2$1$1

.SUBCKT nfet$5$1$2$1$1 \$1 \$2 \$3
.ENDS nfet$5$1$2$1$1

.SUBCKT vias_gen$16$2$1$2$1$1 \$1
.ENDS vias_gen$16$2$1$2$1$1

.SUBCKT vias_gen$17$2$1$2$1$1 \$1
.ENDS vias_gen$17$2$1$2$1$1

.SUBCKT pfet$5$2$1$2$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$2$1$1

.SUBCKT nfet$3$2$1$2$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$2$1$1

.SUBCKT nfet$3$1$1$1$2$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$2$1$1

.SUBCKT vias_gen$16$1$1$1$2$1$1 \$1
.ENDS vias_gen$16$1$1$1$2$1$1

.SUBCKT nfet$4$1$1$2$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$1$2$1$1

.SUBCKT vias_gen$15$1$1$1$2$1$1 \$1
.ENDS vias_gen$15$1$1$1$2$1$1

.SUBCKT vias_gen$14$1$1$1$2$1$1 \$1
.ENDS vias_gen$14$1$1$1$2$1$1

.SUBCKT pfet$4$1$1$1$2$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$2$1$1

.SUBCKT vias_gen$13$1$1$1$2$1$1 \$1
.ENDS vias_gen$13$1$1$1$2$1$1

.SUBCKT vias_gen$12$1$1$1$2$1$1 \$1
.ENDS vias_gen$12$1$1$1$2$1$1

.SUBCKT pfet$5$1$1$1$2$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$2$1$1

.SUBCKT vias_gen$8$1$1$1$2$1$1 \$1
.ENDS vias_gen$8$1$1$1$2$1$1

.SUBCKT vias_gen$17$1$1$1$2$1$1 \$1
.ENDS vias_gen$17$1$1$1$2$1$1

.SUBCKT vias_gen$8$3$2$1$1 \$1
.ENDS vias_gen$8$3$2$1$1

.SUBCKT vias_gen$13$3$2$1$1 \$1
.ENDS vias_gen$13$3$2$1$1

.SUBCKT vias_gen$12$3$2$1$1 \$1
.ENDS vias_gen$12$3$2$1$1

.SUBCKT vias_gen$14$3$2$1$1 \$1
.ENDS vias_gen$14$3$2$1$1

.SUBCKT pfet$4$3$2$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$2$1$1

.SUBCKT vias_gen$15$3$2$1$1 \$1
.ENDS vias_gen$15$3$2$1$1

.SUBCKT nfet$6$2$1$1 \$1 \$2 \$3
.ENDS nfet$6$2$1$1

.SUBCKT vias_gen$16$3$2$1$1 \$1
.ENDS vias_gen$16$3$2$1$1

.SUBCKT vias_gen$17$3$2$1$1 \$1
.ENDS vias_gen$17$3$2$1$1

.SUBCKT pfet$5$3$2$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$2$1$1

.SUBCKT nfet$3$3$2$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$2$1$1

.SUBCKT nfet$3$1$2$2$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$2$1$1

.SUBCKT vias_gen$16$1$2$2$1$1 \$1
.ENDS vias_gen$16$1$2$2$1$1

.SUBCKT nfet$4$2$2$1$1 \$1 \$2 \$3
.ENDS nfet$4$2$2$1$1

.SUBCKT vias_gen$15$1$2$2$1$1 \$1
.ENDS vias_gen$15$1$2$2$1$1

.SUBCKT vias_gen$14$1$2$2$1$1 \$1
.ENDS vias_gen$14$1$2$2$1$1

.SUBCKT pfet$4$1$2$2$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$2$1$1

.SUBCKT vias_gen$13$1$2$2$1$1 \$1
.ENDS vias_gen$13$1$2$2$1$1

.SUBCKT vias_gen$12$1$2$2$1$1 \$1
.ENDS vias_gen$12$1$2$2$1$1

.SUBCKT pfet$5$1$2$2$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$2$1$1

.SUBCKT vias_gen$8$1$2$2$1$1 \$1
.ENDS vias_gen$8$1$2$2$1$1

.SUBCKT vias_gen$17$1$2$2$1$1 \$1
.ENDS vias_gen$17$1$2$2$1$1

.SUBCKT vias_gen$8$2$1$1$1$2 \$1
.ENDS vias_gen$8$2$1$1$1$2

.SUBCKT vias_gen$13$2$1$1$1$2 \$1
.ENDS vias_gen$13$2$1$1$1$2

.SUBCKT vias_gen$12$2$1$1$1$2 \$1
.ENDS vias_gen$12$2$1$1$1$2

.SUBCKT vias_gen$14$2$1$1$1$2 \$1
.ENDS vias_gen$14$2$1$1$1$2

.SUBCKT pfet$4$2$1$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$1$1$2

.SUBCKT vias_gen$15$2$1$1$1$2 \$1
.ENDS vias_gen$15$2$1$1$1$2

.SUBCKT nfet$5$1$1$1$2 \$1 \$2 \$3
.ENDS nfet$5$1$1$1$2

.SUBCKT vias_gen$16$2$1$1$1$2 \$1
.ENDS vias_gen$16$2$1$1$1$2

.SUBCKT vias_gen$17$2$1$1$1$2 \$1
.ENDS vias_gen$17$2$1$1$1$2

.SUBCKT pfet$5$2$1$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$1$1$2

.SUBCKT nfet$3$2$1$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$1$1$2

.SUBCKT nfet$3$1$1$1$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$1$1$2

.SUBCKT vias_gen$16$1$1$1$1$1$2 \$1
.ENDS vias_gen$16$1$1$1$1$1$2

.SUBCKT nfet$4$1$1$1$1$2 \$1 \$2 \$3
.ENDS nfet$4$1$1$1$1$2

.SUBCKT vias_gen$15$1$1$1$1$1$2 \$1
.ENDS vias_gen$15$1$1$1$1$1$2

.SUBCKT vias_gen$14$1$1$1$1$1$2 \$1
.ENDS vias_gen$14$1$1$1$1$1$2

.SUBCKT pfet$4$1$1$1$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$1$1$2

.SUBCKT vias_gen$13$1$1$1$1$1$2 \$1
.ENDS vias_gen$13$1$1$1$1$1$2

.SUBCKT vias_gen$12$1$1$1$1$1$2 \$1
.ENDS vias_gen$12$1$1$1$1$1$2

.SUBCKT pfet$5$1$1$1$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$1$1$2

.SUBCKT vias_gen$8$1$1$1$1$1$2 \$1
.ENDS vias_gen$8$1$1$1$1$1$2

.SUBCKT vias_gen$17$1$1$1$1$1$2 \$1
.ENDS vias_gen$17$1$1$1$1$1$2

.SUBCKT vias_gen$8$3$1$1$2 \$1
.ENDS vias_gen$8$3$1$1$2

.SUBCKT vias_gen$13$3$1$1$2 \$1
.ENDS vias_gen$13$3$1$1$2

.SUBCKT vias_gen$12$3$1$1$2 \$1
.ENDS vias_gen$12$3$1$1$2

.SUBCKT vias_gen$14$3$1$1$2 \$1
.ENDS vias_gen$14$3$1$1$2

.SUBCKT pfet$4$3$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$1$1$2

.SUBCKT vias_gen$15$3$1$1$2 \$1
.ENDS vias_gen$15$3$1$1$2

.SUBCKT nfet$6$1$1$2 \$1 \$2 \$3
.ENDS nfet$6$1$1$2

.SUBCKT vias_gen$16$3$1$1$2 \$1
.ENDS vias_gen$16$3$1$1$2

.SUBCKT vias_gen$17$3$1$1$2 \$1
.ENDS vias_gen$17$3$1$1$2

.SUBCKT pfet$5$3$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$1$1$2

.SUBCKT nfet$3$3$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$1$1$2

.SUBCKT nfet$3$1$2$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$1$1$2

.SUBCKT vias_gen$16$1$2$1$1$2 \$1
.ENDS vias_gen$16$1$2$1$1$2

.SUBCKT nfet$4$2$1$1$2 \$1 \$2 \$3
.ENDS nfet$4$2$1$1$2

.SUBCKT vias_gen$15$1$2$1$1$2 \$1
.ENDS vias_gen$15$1$2$1$1$2

.SUBCKT vias_gen$14$1$2$1$1$2 \$1
.ENDS vias_gen$14$1$2$1$1$2

.SUBCKT pfet$4$1$2$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$1$1$2

.SUBCKT vias_gen$13$1$2$1$1$2 \$1
.ENDS vias_gen$13$1$2$1$1$2

.SUBCKT vias_gen$12$1$2$1$1$2 \$1
.ENDS vias_gen$12$1$2$1$1$2

.SUBCKT pfet$5$1$2$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$1$1$2

.SUBCKT vias_gen$8$1$2$1$1$2 \$1
.ENDS vias_gen$8$1$2$1$1$2

.SUBCKT vias_gen$17$1$2$1$1$2 \$1
.ENDS vias_gen$17$1$2$1$1$2

.SUBCKT vias_gen$8$2$2$1$2 \$1
.ENDS vias_gen$8$2$2$1$2

.SUBCKT vias_gen$13$2$2$1$2 \$1
.ENDS vias_gen$13$2$2$1$2

.SUBCKT vias_gen$12$2$2$1$2 \$1
.ENDS vias_gen$12$2$2$1$2

.SUBCKT vias_gen$14$2$2$1$2 \$1
.ENDS vias_gen$14$2$2$1$2

.SUBCKT pfet$4$2$2$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$2$1$2

.SUBCKT vias_gen$15$2$2$1$2 \$1
.ENDS vias_gen$15$2$2$1$2

.SUBCKT nfet$5$2$1$2 \$1 \$2 \$3
.ENDS nfet$5$2$1$2

.SUBCKT vias_gen$16$2$2$1$2 \$1
.ENDS vias_gen$16$2$2$1$2

.SUBCKT vias_gen$17$2$2$1$2 \$1
.ENDS vias_gen$17$2$2$1$2

.SUBCKT pfet$5$2$2$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$2$1$2

.SUBCKT nfet$3$2$2$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$2$1$2

.SUBCKT nfet$3$1$1$2$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$2$1$2

.SUBCKT vias_gen$16$1$1$2$1$2 \$1
.ENDS vias_gen$16$1$1$2$1$2

.SUBCKT nfet$4$1$2$1$2 \$1 \$2 \$3
.ENDS nfet$4$1$2$1$2

.SUBCKT vias_gen$15$1$1$2$1$2 \$1
.ENDS vias_gen$15$1$1$2$1$2

.SUBCKT vias_gen$14$1$1$2$1$2 \$1
.ENDS vias_gen$14$1$1$2$1$2

.SUBCKT pfet$4$1$1$2$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$2$1$2

.SUBCKT vias_gen$13$1$1$2$1$2 \$1
.ENDS vias_gen$13$1$1$2$1$2

.SUBCKT vias_gen$12$1$1$2$1$2 \$1
.ENDS vias_gen$12$1$1$2$1$2

.SUBCKT pfet$5$1$1$2$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$2$1$2

.SUBCKT vias_gen$8$1$1$2$1$2 \$1
.ENDS vias_gen$8$1$1$2$1$2

.SUBCKT vias_gen$17$1$1$2$1$2 \$1
.ENDS vias_gen$17$1$1$2$1$2

.SUBCKT vias_gen$8$2$1$2$2 \$1
.ENDS vias_gen$8$2$1$2$2

.SUBCKT vias_gen$13$2$1$2$2 \$1
.ENDS vias_gen$13$2$1$2$2

.SUBCKT vias_gen$12$2$1$2$2 \$1
.ENDS vias_gen$12$2$1$2$2

.SUBCKT vias_gen$14$2$1$2$2 \$1
.ENDS vias_gen$14$2$1$2$2

.SUBCKT pfet$4$2$1$2$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$2$2

.SUBCKT vias_gen$15$2$1$2$2 \$1
.ENDS vias_gen$15$2$1$2$2

.SUBCKT nfet$5$1$2$2 \$1 \$2 \$3
.ENDS nfet$5$1$2$2

.SUBCKT vias_gen$16$2$1$2$2 \$1
.ENDS vias_gen$16$2$1$2$2

.SUBCKT vias_gen$17$2$1$2$2 \$1
.ENDS vias_gen$17$2$1$2$2

.SUBCKT pfet$5$2$1$2$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$2$2

.SUBCKT nfet$3$2$1$2$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$2$2

.SUBCKT nfet$3$1$1$1$2$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$2$2

.SUBCKT vias_gen$16$1$1$1$2$2 \$1
.ENDS vias_gen$16$1$1$1$2$2

.SUBCKT nfet$4$1$1$2$2 \$1 \$2 \$3
.ENDS nfet$4$1$1$2$2

.SUBCKT vias_gen$15$1$1$1$2$2 \$1
.ENDS vias_gen$15$1$1$1$2$2

.SUBCKT vias_gen$14$1$1$1$2$2 \$1
.ENDS vias_gen$14$1$1$1$2$2

.SUBCKT pfet$4$1$1$1$2$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$2$2

.SUBCKT vias_gen$13$1$1$1$2$2 \$1
.ENDS vias_gen$13$1$1$1$2$2

.SUBCKT vias_gen$12$1$1$1$2$2 \$1
.ENDS vias_gen$12$1$1$1$2$2

.SUBCKT pfet$5$1$1$1$2$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$2$2

.SUBCKT vias_gen$8$1$1$1$2$2 \$1
.ENDS vias_gen$8$1$1$1$2$2

.SUBCKT vias_gen$17$1$1$1$2$2 \$1
.ENDS vias_gen$17$1$1$1$2$2

.SUBCKT vias_gen$8$3$2$2 \$1
.ENDS vias_gen$8$3$2$2

.SUBCKT vias_gen$13$3$2$2 \$1
.ENDS vias_gen$13$3$2$2

.SUBCKT vias_gen$12$3$2$2 \$1
.ENDS vias_gen$12$3$2$2

.SUBCKT vias_gen$14$3$2$2 \$1
.ENDS vias_gen$14$3$2$2

.SUBCKT pfet$4$3$2$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$2$2

.SUBCKT vias_gen$15$3$2$2 \$1
.ENDS vias_gen$15$3$2$2

.SUBCKT nfet$6$2$2 \$1 \$2 \$3
.ENDS nfet$6$2$2

.SUBCKT vias_gen$16$3$2$2 \$1
.ENDS vias_gen$16$3$2$2

.SUBCKT vias_gen$17$3$2$2 \$1
.ENDS vias_gen$17$3$2$2

.SUBCKT pfet$5$3$2$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$2$2

.SUBCKT nfet$3$3$2$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$2$2

.SUBCKT nfet$3$1$2$2$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$2$2

.SUBCKT vias_gen$16$1$2$2$2 \$1
.ENDS vias_gen$16$1$2$2$2

.SUBCKT nfet$4$2$2$2 \$1 \$2 \$3
.ENDS nfet$4$2$2$2

.SUBCKT vias_gen$15$1$2$2$2 \$1
.ENDS vias_gen$15$1$2$2$2

.SUBCKT vias_gen$14$1$2$2$2 \$1
.ENDS vias_gen$14$1$2$2$2

.SUBCKT pfet$4$1$2$2$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$2$2

.SUBCKT vias_gen$13$1$2$2$2 \$1
.ENDS vias_gen$13$1$2$2$2

.SUBCKT vias_gen$12$1$2$2$2 \$1
.ENDS vias_gen$12$1$2$2$2

.SUBCKT pfet$5$1$2$2$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$2$2

.SUBCKT vias_gen$8$1$2$2$2 \$1
.ENDS vias_gen$8$1$2$2$2

.SUBCKT vias_gen$17$1$2$2$2 \$1
.ENDS vias_gen$17$1$2$2$2

.SUBCKT vias_gen$8$3$1$1$1 \$1
.ENDS vias_gen$8$3$1$1$1

.SUBCKT vias_gen$13$3$1$1$1 \$1
.ENDS vias_gen$13$3$1$1$1

.SUBCKT vias_gen$12$3$1$1$1 \$1
.ENDS vias_gen$12$3$1$1$1

.SUBCKT vias_gen$14$3$1$1$1 \$1
.ENDS vias_gen$14$3$1$1$1

.SUBCKT pfet$4$3$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$1$1$1

.SUBCKT vias_gen$15$3$1$1$1 \$1
.ENDS vias_gen$15$3$1$1$1

.SUBCKT nfet$6$1$1$1 \$1 \$2 \$3
.ENDS nfet$6$1$1$1

.SUBCKT vias_gen$16$3$1$1$1 \$1
.ENDS vias_gen$16$3$1$1$1

.SUBCKT vias_gen$17$3$1$1$1 \$1
.ENDS vias_gen$17$3$1$1$1

.SUBCKT pfet$5$3$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$1$1$1

.SUBCKT nfet$3$3$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$1$1$1

.SUBCKT nfet$3$1$2$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$1$1$1

.SUBCKT vias_gen$16$1$2$1$1$1 \$1
.ENDS vias_gen$16$1$2$1$1$1

.SUBCKT nfet$4$2$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$2$1$1$1

.SUBCKT vias_gen$15$1$2$1$1$1 \$1
.ENDS vias_gen$15$1$2$1$1$1

.SUBCKT vias_gen$14$1$2$1$1$1 \$1
.ENDS vias_gen$14$1$2$1$1$1

.SUBCKT pfet$4$1$2$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$1$1$1

.SUBCKT vias_gen$13$1$2$1$1$1 \$1
.ENDS vias_gen$13$1$2$1$1$1

.SUBCKT vias_gen$12$1$2$1$1$1 \$1
.ENDS vias_gen$12$1$2$1$1$1

.SUBCKT pfet$5$1$2$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$1$1$1

.SUBCKT vias_gen$8$1$2$1$1$1 \$1
.ENDS vias_gen$8$1$2$1$1$1

.SUBCKT vias_gen$17$1$2$1$1$1 \$1
.ENDS vias_gen$17$1$2$1$1$1

.SUBCKT vias_gen$8$2$2$1$1 \$1
.ENDS vias_gen$8$2$2$1$1

.SUBCKT vias_gen$13$2$2$1$1 \$1
.ENDS vias_gen$13$2$2$1$1

.SUBCKT vias_gen$12$2$2$1$1 \$1
.ENDS vias_gen$12$2$2$1$1

.SUBCKT vias_gen$14$2$2$1$1 \$1
.ENDS vias_gen$14$2$2$1$1

.SUBCKT pfet$4$2$2$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$2$1$1

.SUBCKT vias_gen$15$2$2$1$1 \$1
.ENDS vias_gen$15$2$2$1$1

.SUBCKT nfet$5$2$1$1 \$1 \$2 \$3
.ENDS nfet$5$2$1$1

.SUBCKT vias_gen$16$2$2$1$1 \$1
.ENDS vias_gen$16$2$2$1$1

.SUBCKT vias_gen$17$2$2$1$1 \$1
.ENDS vias_gen$17$2$2$1$1

.SUBCKT pfet$5$2$2$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$2$1$1

.SUBCKT nfet$3$2$2$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$2$1$1

.SUBCKT nfet$3$1$1$2$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$2$1$1

.SUBCKT vias_gen$16$1$1$2$1$1 \$1
.ENDS vias_gen$16$1$1$2$1$1

.SUBCKT nfet$4$1$2$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$2$1$1

.SUBCKT vias_gen$15$1$1$2$1$1 \$1
.ENDS vias_gen$15$1$1$2$1$1

.SUBCKT vias_gen$14$1$1$2$1$1 \$1
.ENDS vias_gen$14$1$1$2$1$1

.SUBCKT pfet$4$1$1$2$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$2$1$1

.SUBCKT vias_gen$13$1$1$2$1$1 \$1
.ENDS vias_gen$13$1$1$2$1$1

.SUBCKT vias_gen$12$1$1$2$1$1 \$1
.ENDS vias_gen$12$1$1$2$1$1

.SUBCKT pfet$5$1$1$2$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$2$1$1

.SUBCKT vias_gen$8$1$1$2$1$1 \$1
.ENDS vias_gen$8$1$1$2$1$1

.SUBCKT vias_gen$17$1$1$2$1$1 \$1
.ENDS vias_gen$17$1$1$2$1$1

.SUBCKT vias_gen$8$2$1$2$1 \$1
.ENDS vias_gen$8$2$1$2$1

.SUBCKT vias_gen$13$2$1$2$1 \$1
.ENDS vias_gen$13$2$1$2$1

.SUBCKT vias_gen$12$2$1$2$1 \$1
.ENDS vias_gen$12$2$1$2$1

.SUBCKT vias_gen$14$2$1$2$1 \$1
.ENDS vias_gen$14$2$1$2$1

.SUBCKT pfet$4$2$1$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$2$1

.SUBCKT vias_gen$15$2$1$2$1 \$1
.ENDS vias_gen$15$2$1$2$1

.SUBCKT nfet$5$1$2$1 \$1 \$2 \$3
.ENDS nfet$5$1$2$1

.SUBCKT vias_gen$16$2$1$2$1 \$1
.ENDS vias_gen$16$2$1$2$1

.SUBCKT vias_gen$17$2$1$2$1 \$1
.ENDS vias_gen$17$2$1$2$1

.SUBCKT pfet$5$2$1$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$2$1

.SUBCKT nfet$3$2$1$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$2$1

.SUBCKT nfet$3$1$1$1$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$2$1

.SUBCKT vias_gen$16$1$1$1$2$1 \$1
.ENDS vias_gen$16$1$1$1$2$1

.SUBCKT nfet$4$1$1$2$1 \$1 \$2 \$3
.ENDS nfet$4$1$1$2$1

.SUBCKT vias_gen$15$1$1$1$2$1 \$1
.ENDS vias_gen$15$1$1$1$2$1

.SUBCKT vias_gen$14$1$1$1$2$1 \$1
.ENDS vias_gen$14$1$1$1$2$1

.SUBCKT pfet$4$1$1$1$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$2$1

.SUBCKT vias_gen$13$1$1$1$2$1 \$1
.ENDS vias_gen$13$1$1$1$2$1

.SUBCKT vias_gen$12$1$1$1$2$1 \$1
.ENDS vias_gen$12$1$1$1$2$1

.SUBCKT pfet$5$1$1$1$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$2$1

.SUBCKT vias_gen$8$1$1$1$2$1 \$1
.ENDS vias_gen$8$1$1$1$2$1

.SUBCKT vias_gen$17$1$1$1$2$1 \$1
.ENDS vias_gen$17$1$1$1$2$1

.SUBCKT vias_gen$8$3$2$1 \$1
.ENDS vias_gen$8$3$2$1

.SUBCKT vias_gen$13$3$2$1 \$1
.ENDS vias_gen$13$3$2$1

.SUBCKT vias_gen$12$3$2$1 \$1
.ENDS vias_gen$12$3$2$1

.SUBCKT vias_gen$14$3$2$1 \$1
.ENDS vias_gen$14$3$2$1

.SUBCKT pfet$4$3$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$2$1

.SUBCKT vias_gen$15$3$2$1 \$1
.ENDS vias_gen$15$3$2$1

.SUBCKT nfet$6$2$1 \$1 \$2 \$3
.ENDS nfet$6$2$1

.SUBCKT vias_gen$16$3$2$1 \$1
.ENDS vias_gen$16$3$2$1

.SUBCKT vias_gen$17$3$2$1 \$1
.ENDS vias_gen$17$3$2$1

.SUBCKT pfet$5$3$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$2$1

.SUBCKT nfet$3$3$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$2$1

.SUBCKT nfet$3$1$2$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$2$1

.SUBCKT vias_gen$16$1$2$2$1 \$1
.ENDS vias_gen$16$1$2$2$1

.SUBCKT nfet$4$2$2$1 \$1 \$2 \$3
.ENDS nfet$4$2$2$1

.SUBCKT vias_gen$15$1$2$2$1 \$1
.ENDS vias_gen$15$1$2$2$1

.SUBCKT vias_gen$14$1$2$2$1 \$1
.ENDS vias_gen$14$1$2$2$1

.SUBCKT pfet$4$1$2$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$2$1

.SUBCKT vias_gen$13$1$2$2$1 \$1
.ENDS vias_gen$13$1$2$2$1

.SUBCKT vias_gen$12$1$2$2$1 \$1
.ENDS vias_gen$12$1$2$2$1

.SUBCKT pfet$5$1$2$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$2$1

.SUBCKT vias_gen$8$1$2$2$1 \$1
.ENDS vias_gen$8$1$2$2$1

.SUBCKT vias_gen$17$1$2$2$1 \$1
.ENDS vias_gen$17$1$2$2$1

.SUBCKT vias_gen$8$2$1$1$1 \$1
.ENDS vias_gen$8$2$1$1$1

.SUBCKT vias_gen$13$2$1$1$1 \$1
.ENDS vias_gen$13$2$1$1$1

.SUBCKT vias_gen$12$2$1$1$1 \$1
.ENDS vias_gen$12$2$1$1$1

.SUBCKT vias_gen$14$2$1$1$1 \$1
.ENDS vias_gen$14$2$1$1$1

.SUBCKT pfet$4$2$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$1$1

.SUBCKT vias_gen$15$2$1$1$1 \$1
.ENDS vias_gen$15$2$1$1$1

.SUBCKT nfet$5$1$1$1 \$1 \$2 \$3
.ENDS nfet$5$1$1$1

.SUBCKT vias_gen$16$2$1$1$1 \$1
.ENDS vias_gen$16$2$1$1$1

.SUBCKT vias_gen$17$2$1$1$1 \$1
.ENDS vias_gen$17$2$1$1$1

.SUBCKT pfet$5$2$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$1$1

.SUBCKT nfet$3$2$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$1$1

.SUBCKT nfet$3$1$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$1$1

.SUBCKT vias_gen$16$1$1$1$1$1 \$1
.ENDS vias_gen$16$1$1$1$1$1

.SUBCKT nfet$4$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$1$1$1

.SUBCKT vias_gen$15$1$1$1$1$1 \$1
.ENDS vias_gen$15$1$1$1$1$1

.SUBCKT vias_gen$14$1$1$1$1$1 \$1
.ENDS vias_gen$14$1$1$1$1$1

.SUBCKT pfet$4$1$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$1$1

.SUBCKT vias_gen$13$1$1$1$1$1 \$1
.ENDS vias_gen$13$1$1$1$1$1

.SUBCKT vias_gen$12$1$1$1$1$1 \$1
.ENDS vias_gen$12$1$1$1$1$1

.SUBCKT pfet$5$1$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$1$1

.SUBCKT vias_gen$8$1$1$1$1$1 \$1
.ENDS vias_gen$8$1$1$1$1$1

.SUBCKT vias_gen$17$1$1$1$1$1 \$1
.ENDS vias_gen$17$1$1$1$1$1

.SUBCKT vias_gen$8$3$1$1 \$1
.ENDS vias_gen$8$3$1$1

.SUBCKT vias_gen$13$3$1$1 \$1
.ENDS vias_gen$13$3$1$1

.SUBCKT vias_gen$12$3$1$1 \$1
.ENDS vias_gen$12$3$1$1

.SUBCKT vias_gen$14$3$1$1 \$1
.ENDS vias_gen$14$3$1$1

.SUBCKT pfet$4$3$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$1$1

.SUBCKT vias_gen$15$3$1$1 \$1
.ENDS vias_gen$15$3$1$1

.SUBCKT nfet$6$1$1 \$1 \$2 \$3
.ENDS nfet$6$1$1

.SUBCKT vias_gen$16$3$1$1 \$1
.ENDS vias_gen$16$3$1$1

.SUBCKT vias_gen$17$3$1$1 \$1
.ENDS vias_gen$17$3$1$1

.SUBCKT pfet$5$3$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$1$1

.SUBCKT nfet$3$3$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$1$1

.SUBCKT nfet$3$1$2$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$1$1

.SUBCKT vias_gen$16$1$2$1$1 \$1
.ENDS vias_gen$16$1$2$1$1

.SUBCKT nfet$4$2$1$1 \$1 \$2 \$3
.ENDS nfet$4$2$1$1

.SUBCKT vias_gen$15$1$2$1$1 \$1
.ENDS vias_gen$15$1$2$1$1

.SUBCKT vias_gen$14$1$2$1$1 \$1
.ENDS vias_gen$14$1$2$1$1

.SUBCKT pfet$4$1$2$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$1$1

.SUBCKT vias_gen$13$1$2$1$1 \$1
.ENDS vias_gen$13$1$2$1$1

.SUBCKT vias_gen$12$1$2$1$1 \$1
.ENDS vias_gen$12$1$2$1$1

.SUBCKT pfet$5$1$2$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$1$1

.SUBCKT vias_gen$8$1$2$1$1 \$1
.ENDS vias_gen$8$1$2$1$1

.SUBCKT vias_gen$17$1$2$1$1 \$1
.ENDS vias_gen$17$1$2$1$1

.SUBCKT vias_gen$8$2$2$1 \$1
.ENDS vias_gen$8$2$2$1

.SUBCKT vias_gen$13$2$2$1 \$1
.ENDS vias_gen$13$2$2$1

.SUBCKT vias_gen$12$2$2$1 \$1
.ENDS vias_gen$12$2$2$1

.SUBCKT vias_gen$14$2$2$1 \$1
.ENDS vias_gen$14$2$2$1

.SUBCKT pfet$4$2$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$2$1

.SUBCKT vias_gen$15$2$2$1 \$1
.ENDS vias_gen$15$2$2$1

.SUBCKT nfet$5$2$1 \$1 \$2 \$3
.ENDS nfet$5$2$1

.SUBCKT vias_gen$16$2$2$1 \$1
.ENDS vias_gen$16$2$2$1

.SUBCKT vias_gen$17$2$2$1 \$1
.ENDS vias_gen$17$2$2$1

.SUBCKT pfet$5$2$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$2$1

.SUBCKT nfet$3$2$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$2$1

.SUBCKT nfet$3$1$1$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$2$1

.SUBCKT vias_gen$16$1$1$2$1 \$1
.ENDS vias_gen$16$1$1$2$1

.SUBCKT nfet$4$1$2$1 \$1 \$2 \$3
.ENDS nfet$4$1$2$1

.SUBCKT vias_gen$15$1$1$2$1 \$1
.ENDS vias_gen$15$1$1$2$1

.SUBCKT vias_gen$14$1$1$2$1 \$1
.ENDS vias_gen$14$1$1$2$1

.SUBCKT pfet$4$1$1$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$2$1

.SUBCKT vias_gen$13$1$1$2$1 \$1
.ENDS vias_gen$13$1$1$2$1

.SUBCKT vias_gen$12$1$1$2$1 \$1
.ENDS vias_gen$12$1$1$2$1

.SUBCKT pfet$5$1$1$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$2$1

.SUBCKT vias_gen$8$1$1$2$1 \$1
.ENDS vias_gen$8$1$1$2$1

.SUBCKT vias_gen$17$1$1$2$1 \$1
.ENDS vias_gen$17$1$1$2$1

.SUBCKT vias_gen$8$2$1$2 \$1
.ENDS vias_gen$8$2$1$2

.SUBCKT vias_gen$13$2$1$2 \$1
.ENDS vias_gen$13$2$1$2

.SUBCKT vias_gen$12$2$1$2 \$1
.ENDS vias_gen$12$2$1$2

.SUBCKT vias_gen$14$2$1$2 \$1
.ENDS vias_gen$14$2$1$2

.SUBCKT pfet$4$2$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$2

.SUBCKT vias_gen$15$2$1$2 \$1
.ENDS vias_gen$15$2$1$2

.SUBCKT nfet$5$1$2 \$1 \$2 \$3
.ENDS nfet$5$1$2

.SUBCKT vias_gen$16$2$1$2 \$1
.ENDS vias_gen$16$2$1$2

.SUBCKT vias_gen$17$2$1$2 \$1
.ENDS vias_gen$17$2$1$2

.SUBCKT pfet$5$2$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$2

.SUBCKT nfet$3$2$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$2

.SUBCKT nfet$3$1$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$2

.SUBCKT vias_gen$16$1$1$1$2 \$1
.ENDS vias_gen$16$1$1$1$2

.SUBCKT nfet$4$1$1$2 \$1 \$2 \$3
.ENDS nfet$4$1$1$2

.SUBCKT vias_gen$15$1$1$1$2 \$1
.ENDS vias_gen$15$1$1$1$2

.SUBCKT vias_gen$14$1$1$1$2 \$1
.ENDS vias_gen$14$1$1$1$2

.SUBCKT pfet$4$1$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$2

.SUBCKT vias_gen$13$1$1$1$2 \$1
.ENDS vias_gen$13$1$1$1$2

.SUBCKT vias_gen$12$1$1$1$2 \$1
.ENDS vias_gen$12$1$1$1$2

.SUBCKT pfet$5$1$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$2

.SUBCKT vias_gen$8$1$1$1$2 \$1
.ENDS vias_gen$8$1$1$1$2

.SUBCKT vias_gen$17$1$1$1$2 \$1
.ENDS vias_gen$17$1$1$1$2

.SUBCKT vias_gen$8$3$2 \$1
.ENDS vias_gen$8$3$2

.SUBCKT vias_gen$13$3$2 \$1
.ENDS vias_gen$13$3$2

.SUBCKT vias_gen$12$3$2 \$1
.ENDS vias_gen$12$3$2

.SUBCKT vias_gen$14$3$2 \$1
.ENDS vias_gen$14$3$2

.SUBCKT pfet$4$3$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$2

.SUBCKT vias_gen$15$3$2 \$1
.ENDS vias_gen$15$3$2

.SUBCKT nfet$6$2 \$1 \$2 \$3
.ENDS nfet$6$2

.SUBCKT vias_gen$16$3$2 \$1
.ENDS vias_gen$16$3$2

.SUBCKT vias_gen$17$3$2 \$1
.ENDS vias_gen$17$3$2

.SUBCKT pfet$5$3$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$2

.SUBCKT nfet$3$3$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$2

.SUBCKT nfet$3$1$2$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$2

.SUBCKT vias_gen$16$1$2$2 \$1
.ENDS vias_gen$16$1$2$2

.SUBCKT nfet$4$2$2 \$1 \$2 \$3
.ENDS nfet$4$2$2

.SUBCKT vias_gen$15$1$2$2 \$1
.ENDS vias_gen$15$1$2$2

.SUBCKT vias_gen$14$1$2$2 \$1
.ENDS vias_gen$14$1$2$2

.SUBCKT pfet$4$1$2$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$2

.SUBCKT vias_gen$13$1$2$2 \$1
.ENDS vias_gen$13$1$2$2

.SUBCKT vias_gen$12$1$2$2 \$1
.ENDS vias_gen$12$1$2$2

.SUBCKT pfet$5$1$2$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$2

.SUBCKT vias_gen$8$1$2$2 \$1
.ENDS vias_gen$8$1$2$2

.SUBCKT vias_gen$17$1$2$2 \$1
.ENDS vias_gen$17$1$2$2

.SUBCKT vias_gen$8$2$1$1 \$1
.ENDS vias_gen$8$2$1$1

.SUBCKT vias_gen$13$2$1$1 \$1
.ENDS vias_gen$13$2$1$1

.SUBCKT vias_gen$12$2$1$1 \$1
.ENDS vias_gen$12$2$1$1

.SUBCKT vias_gen$14$2$1$1 \$1
.ENDS vias_gen$14$2$1$1

.SUBCKT pfet$4$2$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$1

.SUBCKT vias_gen$15$2$1$1 \$1
.ENDS vias_gen$15$2$1$1

.SUBCKT nfet$5$1$1 \$1 \$2 \$3
.ENDS nfet$5$1$1

.SUBCKT vias_gen$16$2$1$1 \$1
.ENDS vias_gen$16$2$1$1

.SUBCKT vias_gen$17$2$1$1 \$1
.ENDS vias_gen$17$2$1$1

.SUBCKT pfet$5$2$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$1

.SUBCKT nfet$3$2$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$1

.SUBCKT nfet$3$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$1

.SUBCKT vias_gen$16$1$1$1$1 \$1
.ENDS vias_gen$16$1$1$1$1

.SUBCKT nfet$4$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$1$1

.SUBCKT vias_gen$15$1$1$1$1 \$1
.ENDS vias_gen$15$1$1$1$1

.SUBCKT vias_gen$14$1$1$1$1 \$1
.ENDS vias_gen$14$1$1$1$1

.SUBCKT pfet$4$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$1

.SUBCKT vias_gen$13$1$1$1$1 \$1
.ENDS vias_gen$13$1$1$1$1

.SUBCKT vias_gen$12$1$1$1$1 \$1
.ENDS vias_gen$12$1$1$1$1

.SUBCKT pfet$5$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$1

.SUBCKT vias_gen$8$1$1$1$1 \$1
.ENDS vias_gen$8$1$1$1$1

.SUBCKT vias_gen$17$1$1$1$1 \$1
.ENDS vias_gen$17$1$1$1$1

.SUBCKT vias_gen$8$3$1 \$1
.ENDS vias_gen$8$3$1

.SUBCKT vias_gen$13$3$1 \$1
.ENDS vias_gen$13$3$1

.SUBCKT vias_gen$12$3$1 \$1
.ENDS vias_gen$12$3$1

.SUBCKT vias_gen$14$3$1 \$1
.ENDS vias_gen$14$3$1

.SUBCKT pfet$4$3$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$3$1

.SUBCKT vias_gen$15$3$1 \$1
.ENDS vias_gen$15$3$1

.SUBCKT nfet$6$1 \$1 \$2 \$3
.ENDS nfet$6$1

.SUBCKT vias_gen$16$3$1 \$1
.ENDS vias_gen$16$3$1

.SUBCKT vias_gen$17$3$1 \$1
.ENDS vias_gen$17$3$1

.SUBCKT pfet$5$3$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3$1

.SUBCKT nfet$3$3$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3$1

.SUBCKT nfet$3$1$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2$1

.SUBCKT vias_gen$16$1$2$1 \$1
.ENDS vias_gen$16$1$2$1

.SUBCKT nfet$4$2$1 \$1 \$2 \$3
.ENDS nfet$4$2$1

.SUBCKT vias_gen$15$1$2$1 \$1
.ENDS vias_gen$15$1$2$1

.SUBCKT vias_gen$14$1$2$1 \$1
.ENDS vias_gen$14$1$2$1

.SUBCKT pfet$4$1$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2$1

.SUBCKT vias_gen$13$1$2$1 \$1
.ENDS vias_gen$13$1$2$1

.SUBCKT vias_gen$12$1$2$1 \$1
.ENDS vias_gen$12$1$2$1

.SUBCKT pfet$5$1$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2$1

.SUBCKT vias_gen$8$1$2$1 \$1
.ENDS vias_gen$8$1$2$1

.SUBCKT vias_gen$17$1$2$1 \$1
.ENDS vias_gen$17$1$2$1

.SUBCKT vias_gen$8$2$2 \$1
.ENDS vias_gen$8$2$2

.SUBCKT vias_gen$13$2$2 \$1
.ENDS vias_gen$13$2$2

.SUBCKT vias_gen$12$2$2 \$1
.ENDS vias_gen$12$2$2

.SUBCKT vias_gen$14$2$2 \$1
.ENDS vias_gen$14$2$2

.SUBCKT pfet$4$2$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$2

.SUBCKT vias_gen$15$2$2 \$1
.ENDS vias_gen$15$2$2

.SUBCKT nfet$5$2 \$1 \$2 \$3
.ENDS nfet$5$2

.SUBCKT vias_gen$16$2$2 \$1
.ENDS vias_gen$16$2$2

.SUBCKT vias_gen$17$2$2 \$1
.ENDS vias_gen$17$2$2

.SUBCKT pfet$5$2$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$2

.SUBCKT nfet$3$2$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$2

.SUBCKT nfet$3$1$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$2

.SUBCKT vias_gen$16$1$1$2 \$1
.ENDS vias_gen$16$1$1$2

.SUBCKT nfet$4$1$2 \$1 \$2 \$3
.ENDS nfet$4$1$2

.SUBCKT vias_gen$15$1$1$2 \$1
.ENDS vias_gen$15$1$1$2

.SUBCKT vias_gen$14$1$1$2 \$1
.ENDS vias_gen$14$1$1$2

.SUBCKT pfet$4$1$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$2

.SUBCKT vias_gen$13$1$1$2 \$1
.ENDS vias_gen$13$1$1$2

.SUBCKT vias_gen$12$1$1$2 \$1
.ENDS vias_gen$12$1$1$2

.SUBCKT pfet$5$1$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$2

.SUBCKT vias_gen$8$1$1$2 \$1
.ENDS vias_gen$8$1$1$2

.SUBCKT vias_gen$17$1$1$2 \$1
.ENDS vias_gen$17$1$1$2

.SUBCKT vias_gen$8$2$1 \$1
.ENDS vias_gen$8$2$1

.SUBCKT vias_gen$13$2$1 \$1
.ENDS vias_gen$13$2$1

.SUBCKT vias_gen$12$2$1 \$1
.ENDS vias_gen$12$2$1

.SUBCKT vias_gen$14$2$1 \$1
.ENDS vias_gen$14$2$1

.SUBCKT pfet$4$2$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1

.SUBCKT vias_gen$15$2$1 \$1
.ENDS vias_gen$15$2$1

.SUBCKT nfet$5$1 \$1 \$2 \$3
.ENDS nfet$5$1

.SUBCKT vias_gen$16$2$1 \$1
.ENDS vias_gen$16$2$1

.SUBCKT vias_gen$17$2$1 \$1
.ENDS vias_gen$17$2$1

.SUBCKT pfet$5$2$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1

.SUBCKT nfet$3$2$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1

.SUBCKT nfet$3$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1

.SUBCKT vias_gen$16$1$1$1 \$1
.ENDS vias_gen$16$1$1$1

.SUBCKT nfet$4$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$1

.SUBCKT vias_gen$15$1$1$1 \$1
.ENDS vias_gen$15$1$1$1

.SUBCKT vias_gen$14$1$1$1 \$1
.ENDS vias_gen$14$1$1$1

.SUBCKT pfet$4$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1

.SUBCKT vias_gen$13$1$1$1 \$1
.ENDS vias_gen$13$1$1$1

.SUBCKT vias_gen$12$1$1$1 \$1
.ENDS vias_gen$12$1$1$1

.SUBCKT pfet$5$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1

.SUBCKT vias_gen$8$1$1$1 \$1
.ENDS vias_gen$8$1$1$1

.SUBCKT vias_gen$17$1$1$1 \$1
.ENDS vias_gen$17$1$1$1

.SUBCKT vias_gen$8$3 \$1
.ENDS vias_gen$8$3

.SUBCKT vias_gen$13$3 \$1
.ENDS vias_gen$13$3

.SUBCKT vias_gen$12$3 \$1
.ENDS vias_gen$12$3

.SUBCKT vias_gen$14$3 \$1
.ENDS vias_gen$14$3

.SUBCKT pfet$4$3 \$1 \$2 \$3 \$4
.ENDS pfet$4$3

.SUBCKT vias_gen$15$3 \$1
.ENDS vias_gen$15$3

.SUBCKT nfet$6 \$1 \$2 \$3
.ENDS nfet$6

.SUBCKT vias_gen$16$3 \$1
.ENDS vias_gen$16$3

.SUBCKT vias_gen$17$3 \$1
.ENDS vias_gen$17$3

.SUBCKT pfet$5$3 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$3

.SUBCKT nfet$3$3 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$3

.SUBCKT nfet$3$1$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$2

.SUBCKT vias_gen$16$1$2 \$1
.ENDS vias_gen$16$1$2

.SUBCKT nfet$4$2 \$1 \$2 \$3
.ENDS nfet$4$2

.SUBCKT vias_gen$15$1$2 \$1
.ENDS vias_gen$15$1$2

.SUBCKT vias_gen$14$1$2 \$1
.ENDS vias_gen$14$1$2

.SUBCKT pfet$4$1$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$2

.SUBCKT vias_gen$13$1$2 \$1
.ENDS vias_gen$13$1$2

.SUBCKT vias_gen$12$1$2 \$1
.ENDS vias_gen$12$1$2

.SUBCKT pfet$5$1$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$2

.SUBCKT vias_gen$8$1$2 \$1
.ENDS vias_gen$8$1$2

.SUBCKT vias_gen$17$1$2 \$1
.ENDS vias_gen$17$1$2

.SUBCKT vias_gen$8$2 \$1
.ENDS vias_gen$8$2

.SUBCKT vias_gen$13$2 \$1
.ENDS vias_gen$13$2

.SUBCKT vias_gen$12$2 \$1
.ENDS vias_gen$12$2

.SUBCKT vias_gen$14$2 \$1
.ENDS vias_gen$14$2

.SUBCKT pfet$4$2 \$1 \$2 \$3 \$4
.ENDS pfet$4$2

.SUBCKT vias_gen$15$2 \$1
.ENDS vias_gen$15$2

.SUBCKT nfet$5 \$1 \$2 \$3
.ENDS nfet$5

.SUBCKT vias_gen$16$2 \$1
.ENDS vias_gen$16$2

.SUBCKT vias_gen$17$2 \$1
.ENDS vias_gen$17$2

.SUBCKT pfet$5$2 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2

.SUBCKT nfet$3$2 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2

.SUBCKT nfet$3$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1

.SUBCKT vias_gen$16$1$1 \$1
.ENDS vias_gen$16$1$1

.SUBCKT nfet$4$1 \$1 \$2 \$3
.ENDS nfet$4$1

.SUBCKT vias_gen$15$1$1 \$1
.ENDS vias_gen$15$1$1

.SUBCKT vias_gen$14$1$1 \$1
.ENDS vias_gen$14$1$1

.SUBCKT pfet$4$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1

.SUBCKT vias_gen$13$1$1 \$1
.ENDS vias_gen$13$1$1

.SUBCKT vias_gen$12$1$1 \$1
.ENDS vias_gen$12$1$1

.SUBCKT pfet$5$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1

.SUBCKT vias_gen$8$1$1 \$1
.ENDS vias_gen$8$1$1

.SUBCKT vias_gen$17$1$1 \$1
.ENDS vias_gen$17$1$1

.SUBCKT vias_gen$8 \$1
.ENDS vias_gen$8

.SUBCKT vias_gen$13 \$1
.ENDS vias_gen$13

.SUBCKT vias_gen$12 \$1
.ENDS vias_gen$12

.SUBCKT vias_gen$14 \$1
.ENDS vias_gen$14

.SUBCKT pfet$4 \$1 \$2 \$3 \$4
.ENDS pfet$4

.SUBCKT vias_gen$15 \$1
.ENDS vias_gen$15

.SUBCKT nfet \$1 \$2 \$3
.ENDS nfet

.SUBCKT vias_gen$16 \$1
.ENDS vias_gen$16

.SUBCKT vias_gen$17 \$1
.ENDS vias_gen$17

.SUBCKT pfet$5 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5

.SUBCKT nfet$3 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3

.SUBCKT nfet$3$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1

.SUBCKT vias_gen$16$1 \$1
.ENDS vias_gen$16$1

.SUBCKT nfet$4 \$1 \$2 \$3
.ENDS nfet$4

.SUBCKT vias_gen$15$1 \$1
.ENDS vias_gen$15$1

.SUBCKT vias_gen$14$1 \$1
.ENDS vias_gen$14$1

.SUBCKT pfet$4$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1

.SUBCKT vias_gen$13$1 \$1
.ENDS vias_gen$13$1

.SUBCKT vias_gen$12$1 \$1
.ENDS vias_gen$12$1

.SUBCKT pfet$5$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1

.SUBCKT vias_gen$8$1 \$1
.ENDS vias_gen$8$1

.SUBCKT vias_gen$17$1 \$1
.ENDS vias_gen$17$1

.SUBCKT vias_gen$8$2$1$1$1$1 \$1
.ENDS vias_gen$8$2$1$1$1$1

.SUBCKT vias_gen$13$2$1$1$1$1 \$1
.ENDS vias_gen$13$2$1$1$1$1

.SUBCKT vias_gen$12$2$1$1$1$1 \$1
.ENDS vias_gen$12$2$1$1$1$1

.SUBCKT vias_gen$14$2$1$1$1$1 \$1
.ENDS vias_gen$14$2$1$1$1$1

.SUBCKT pfet$4$2$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$2$1$1$1$1

.SUBCKT vias_gen$15$2$1$1$1$1 \$1
.ENDS vias_gen$15$2$1$1$1$1

.SUBCKT nfet$5$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$5$1$1$1$1

.SUBCKT vias_gen$16$2$1$1$1$1 \$1
.ENDS vias_gen$16$2$1$1$1$1

.SUBCKT vias_gen$17$2$1$1$1$1 \$1
.ENDS vias_gen$17$2$1$1$1$1

.SUBCKT pfet$5$2$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$2$1$1$1$1

.SUBCKT nfet$3$2$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$2$1$1$1$1

.SUBCKT nfet$3$1$1$1$1$1$1 \$2 \$3 \$4 \$5 sky130_gnd
M$1 \$5 \$3 \$4 sky130_gnd sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 AS=0.135
+ AD=0.135 PS=1.5 PD=1.5
.ENDS nfet$3$1$1$1$1$1$1

.SUBCKT vias_gen$16$1$1$1$1$1$1 \$1
.ENDS vias_gen$16$1$1$1$1$1$1

.SUBCKT nfet$4$1$1$1$1$1 \$1 \$2 \$3
.ENDS nfet$4$1$1$1$1$1

.SUBCKT vias_gen$15$1$1$1$1$1$1 \$1
.ENDS vias_gen$15$1$1$1$1$1$1

.SUBCKT vias_gen$14$1$1$1$1$1$1 \$1
.ENDS vias_gen$14$1$1$1$1$1$1

.SUBCKT pfet$4$1$1$1$1$1$1 \$1 \$2 \$3 \$4
.ENDS pfet$4$1$1$1$1$1$1

.SUBCKT vias_gen$13$1$1$1$1$1$1 \$1
.ENDS vias_gen$13$1$1$1$1$1$1

.SUBCKT vias_gen$12$1$1$1$1$1$1 \$1
.ENDS vias_gen$12$1$1$1$1$1$1

.SUBCKT pfet$5$1$1$1$1$1$1 \$1 \$3 \$4 \$5
M$1 \$5 \$3 \$4 \$1 sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 AS=0.135 AD=0.135
+ PS=1.5 PD=1.5
.ENDS pfet$5$1$1$1$1$1$1

.SUBCKT vias_gen$8$1$1$1$1$1$1 \$1
.ENDS vias_gen$8$1$1$1$1$1$1

.SUBCKT vias_gen$17$1$1$1$1$1$1 \$1
.ENDS vias_gen$17$1$1$1$1$1$1
