** sch_path: /foss/designs/RO_Aging_UNICASS/MOS/nmos_lvt.sch
.subckt nmos_lvt VS VG VD VSS
*.PININFO VS:B VG:B VD:B VSS:B
M1 VD VG VS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends
.end
