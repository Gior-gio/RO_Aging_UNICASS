** sch_path: /foss/designs/xschem_pruebas/inv_prueba.sch
.subckt inv_prueba VDD Out In VSS
*.PININFO Out:B In:B VDD:B VSS:B
XM3 Out In VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 Out In VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
.ends
.end
