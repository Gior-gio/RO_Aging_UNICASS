* Extracted by KLayout with SKY130 LVS runset on : 07/11/2024 00:09

.SUBCKT RO_LVT_13St_x10 RO RON GND DUT_Gate DUT_Header DUT_Footer VDD
+ Drain\x20Force Drain_Sense Out
M$1 \$34 \$24 \$25 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$5 VDD RON \$34 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$45 \$36 \$25 \$19 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$49 VDD DUT_Footer \$36 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$89 \$19 RO Drain_Sense VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$93 \$19 RO Drain\x20Force VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$97 \$38 \$19 \$26 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$101 VDD RON \$38 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$141 \$84 VDD \$24 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$142 \$85 VDD \$24 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$143 VDD \$75 \$24 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$147 \$86 VDD \$75 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$148 \$87 VDD \$75 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$149 VDD \$76 \$75 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$153 \$88 VDD \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$154 \$89 VDD \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$155 VDD \$77 \$76 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$159 \$25 RO DUT_Gate VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$160 \$90 VDD \$77 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$161 \$25 RO \$18 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$162 \$91 VDD \$77 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$163 VDD \$78 \$77 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$167 \$92 VDD \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$168 \$93 VDD \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$169 VDD \$79 \$78 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$173 \$94 VDD \$79 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$174 \$95 VDD \$79 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$175 VDD \$80 \$79 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$179 \$96 VDD \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$180 \$97 VDD \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$181 VDD \$81 \$80 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$185 \$98 VDD \$81 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$186 \$99 VDD \$81 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$187 VDD \$82 \$81 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$191 \$100 VDD \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$192 \$101 VDD \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$193 VDD Out \$82 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$197 \$102 VDD Out VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$198 \$103 VDD Out VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$199 VDD \$26 Out VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$203 \$26 VDD GND VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$204 \$26 VDD \$20 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$205 \$25 \$24 \$6 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$207 \$6 RO GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.26e+13 AD=1.26e+13 PS=96000000 PD=96000000
M$227 \$19 \$25 \$11 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$229 \$11 DUT_Header GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.26e+13 AD=1.26e+13 PS=96000000 PD=96000000
M$249 \$19 RON Drain_Sense GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$251 \$19 RON Drain\x20Force GND sky130_fd_pr__nfet_01v8_lvt L=350000
+ W=4200000 AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$253 \$26 \$19 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$255 \$84 GND \$24 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$256 \$85 GND \$24 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$257 \$24 \$75 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$259 \$86 GND \$75 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$260 \$87 GND \$75 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$261 \$75 \$76 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$263 \$88 GND \$76 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$264 \$89 GND \$76 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$265 \$76 \$77 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$267 \$25 RON DUT_Gate GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$268 \$90 GND \$77 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$269 \$25 RON \$18 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$270 \$91 GND \$77 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$271 \$77 \$78 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$273 \$92 GND \$78 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$274 \$93 GND \$78 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$275 \$78 \$79 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$277 \$94 GND \$79 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$278 \$95 GND \$79 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$279 \$79 \$80 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$281 \$96 GND \$80 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$282 \$97 GND \$80 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$283 \$80 \$81 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$285 \$98 GND \$81 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$286 \$99 GND \$81 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$287 \$81 \$82 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$289 \$100 GND \$82 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$290 \$101 GND \$82 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$291 \$82 Out GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$293 \$102 GND Out GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$294 \$103 GND Out GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$295 Out \$26 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$297 \$26 RON GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$298 \$26 RON \$20 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
.ENDS RO_LVT_13St_x10
