* Extracted by KLayout with SKY130 LVS runset on : 09/11/2024 22:33

.SUBCKT DIV IN GND OUT VDD
M$1 \$113 \$1 \$88 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$2 \$14 IN \$88 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$3 \$89 IN \$90 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$4 \$113 \$1 \$90 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$5 \$114 \$2 \$92 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$6 \$21 \$113 \$92 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$7 \$20 \$113 \$93 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$8 \$114 \$2 \$93 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$9 \$115 \$3 \$94 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$10 \$29 \$114 \$94 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$11 \$28 \$114 \$95 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$12 \$115 \$3 \$95 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$13 \$116 \$4 \$96 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$14 \$37 \$115 \$96 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$15 \$36 \$115 \$97 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$16 \$116 \$4 \$97 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$17 \$117 \$5 \$99 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$18 \$44 \$116 \$99 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$19 \$43 \$116 \$100 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$20 \$117 \$5 \$100 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$21 \$118 \$6 \$101 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$22 \$52 \$117 \$101 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$23 \$51 \$117 \$102 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$24 \$118 \$6 \$102 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$25 \$119 \$7 \$104 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$26 \$59 \$118 \$104 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$27 \$58 \$118 \$105 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$28 \$119 \$7 \$105 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$29 \$120 \$8 \$106 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$30 \$67 \$119 \$106 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$31 \$66 \$119 \$107 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$32 \$120 \$8 \$107 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$33 \$121 \$9 \$108 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$34 \$75 \$120 \$108 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$35 \$74 \$120 \$109 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$36 \$121 \$9 \$109 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$37 OUT \$10 \$111 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$38 \$82 \$121 \$111 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$39 \$81 \$121 \$112 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$40 OUT \$10 \$112 VDD sky130_fd_pr__pfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$41 VDD IN \$1 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000 AS=600000000000
+ AD=600000000000 PS=5200000 PD=5200000
M$43 VDD \$88 \$89 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$45 VDD \$89 \$14 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$47 VDD \$90 \$91 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$49 VDD \$91 \$113 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$51 VDD \$113 \$18 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$53 VDD \$113 \$2 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$55 VDD \$92 \$20 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$57 VDD \$20 \$21 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$59 VDD \$93 \$24 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$61 VDD \$24 \$114 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$63 VDD \$114 \$26 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$65 VDD \$114 \$3 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$67 VDD \$94 \$28 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$69 VDD \$28 \$29 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$71 VDD \$95 \$32 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$73 VDD \$32 \$115 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$75 VDD \$115 \$34 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$77 VDD \$115 \$4 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$79 VDD \$96 \$36 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$81 VDD \$36 \$37 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$83 VDD \$97 \$98 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$85 VDD \$98 \$116 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$87 VDD \$116 \$41 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$89 VDD \$116 \$5 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$91 VDD \$99 \$43 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$93 VDD \$43 \$44 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$95 VDD \$100 \$47 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$97 VDD \$47 \$117 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$99 VDD \$117 \$49 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$101 VDD \$117 \$6 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$103 VDD \$101 \$51 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$105 VDD \$51 \$52 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$107 VDD \$102 \$55 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$109 VDD \$55 \$118 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$111 VDD \$118 \$103 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$113 VDD \$118 \$7 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$115 VDD \$104 \$58 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$117 VDD \$58 \$59 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$119 VDD \$105 \$62 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$121 VDD \$62 \$119 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$123 VDD \$119 \$64 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$125 VDD \$119 \$8 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$127 VDD \$106 \$66 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$129 VDD \$66 \$67 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$131 VDD \$107 \$70 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$133 VDD \$70 \$120 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$135 VDD \$120 \$72 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$137 VDD \$120 \$9 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$139 VDD \$108 \$74 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$141 VDD \$74 \$75 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$143 VDD \$109 \$78 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$145 VDD \$78 \$121 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$147 VDD \$121 \$110 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$149 VDD \$121 \$10 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$151 VDD \$111 \$81 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$153 VDD \$81 \$82 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$155 VDD \$112 \$85 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$157 VDD \$85 OUT VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$159 VDD OUT \$87 VDD sky130_fd_pr__pfet_01v8 L=150000 W=2000000
+ AS=600000000000 AD=600000000000 PS=5200000 PD=5200000
M$161 GND IN \$1 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000 AS=300000000000
+ AD=300000000000 PS=2600000 PD=2600000
M$162 GND \$88 \$89 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$163 GND \$89 \$14 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$164 GND \$90 \$91 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$165 GND \$91 \$113 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$166 GND \$113 \$18 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$167 GND \$113 \$2 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$168 GND \$92 \$20 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$169 GND \$20 \$21 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$170 GND \$93 \$24 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$171 GND \$24 \$114 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$172 GND \$114 \$26 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$173 GND \$114 \$3 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$174 GND \$94 \$28 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$175 GND \$28 \$29 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$176 GND \$95 \$32 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$177 GND \$32 \$115 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$178 GND \$115 \$34 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$179 GND \$115 \$4 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$180 GND \$96 \$36 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$181 GND \$36 \$37 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$182 GND \$97 \$98 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$183 GND \$98 \$116 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$184 GND \$116 \$41 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$185 GND \$116 \$5 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$186 GND \$99 \$43 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$187 GND \$43 \$44 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$188 GND \$100 \$47 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$189 GND \$47 \$117 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$190 GND \$117 \$49 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$191 GND \$117 \$6 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$192 GND \$101 \$51 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$193 GND \$51 \$52 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$194 GND \$102 \$55 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$195 GND \$55 \$118 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$196 GND \$118 \$103 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$197 GND \$118 \$7 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$198 GND \$104 \$58 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$199 GND \$58 \$59 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$200 GND \$105 \$62 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$201 GND \$62 \$119 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$202 GND \$119 \$64 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$203 GND \$119 \$8 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$204 GND \$106 \$66 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$205 GND \$66 \$67 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$206 GND \$107 \$70 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$207 GND \$70 \$120 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$208 GND \$120 \$72 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$209 GND \$120 \$9 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$210 GND \$108 \$74 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$211 GND \$74 \$75 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$212 GND \$109 \$78 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$213 GND \$78 \$121 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$214 GND \$121 \$110 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$215 GND \$121 \$10 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$216 GND \$111 \$81 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$217 GND \$81 \$82 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$218 GND \$112 \$85 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$219 GND \$85 OUT GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$220 GND OUT \$87 GND sky130_fd_pr__nfet_01v8 L=150000 W=1000000
+ AS=300000000000 AD=300000000000 PS=2600000 PD=2600000
M$221 \$113 IN \$88 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$222 \$14 \$1 \$88 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$223 \$89 \$1 \$90 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$224 \$113 IN \$90 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$225 \$114 \$113 \$92 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$226 \$21 \$2 \$92 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$227 \$20 \$2 \$93 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$228 \$114 \$113 \$93 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$229 \$115 \$114 \$94 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$230 \$29 \$3 \$94 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$231 \$28 \$3 \$95 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$232 \$115 \$114 \$95 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$233 \$116 \$115 \$96 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$234 \$37 \$4 \$96 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$235 \$36 \$4 \$97 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$236 \$116 \$115 \$97 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$237 \$117 \$116 \$99 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$238 \$44 \$5 \$99 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$239 \$43 \$5 \$100 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$240 \$117 \$116 \$100 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$241 \$118 \$117 \$101 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$242 \$52 \$6 \$101 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$243 \$51 \$6 \$102 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$244 \$118 \$117 \$102 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$245 \$119 \$118 \$104 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$246 \$59 \$7 \$104 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$247 \$58 \$7 \$105 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$248 \$119 \$118 \$105 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$249 \$120 \$119 \$106 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$250 \$67 \$8 \$106 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$251 \$66 \$8 \$107 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$252 \$120 \$119 \$107 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$253 \$121 \$120 \$108 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$254 \$75 \$9 \$108 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$255 \$74 \$9 \$109 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$256 \$121 \$120 \$109 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$257 OUT \$121 \$111 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$258 \$82 \$10 \$111 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$259 \$81 \$10 \$112 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
M$260 OUT \$121 \$112 GND sky130_fd_pr__nfet_01v8 L=150000 W=650000
+ AS=195000000000 AD=195000000000 PS=1900000 PD=1900000
.ENDS DIV
