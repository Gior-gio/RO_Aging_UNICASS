magic
tech sky130A
magscale 1 2
timestamp 1728607134
<< checkpaint >>
rect -40 -3166 2902 -136
<< error_s >>
rect 1046 -584 1052 -420
rect 1106 -586 1112 -420
rect 1046 -1104 1052 -1030
rect 1106 -1104 1112 -1030
rect 1033 -1373 1091 -1367
rect 1033 -1407 1045 -1373
rect 1033 -1413 1091 -1407
rect 1033 -1681 1091 -1675
rect 1033 -1715 1045 -1681
rect 1033 -1721 1091 -1715
<< locali >>
rect 904 -420 1052 -408
rect 904 -584 916 -420
rect 904 -598 1052 -584
rect 1106 -420 1184 -408
rect 1176 -586 1184 -420
rect 1106 -598 1184 -586
rect 904 -1030 1052 -1018
rect 904 -1104 916 -1030
rect 904 -1116 1052 -1104
rect 1106 -1030 1184 -1018
rect 1176 -1104 1184 -1030
rect 1106 -1116 1184 -1104
<< viali >>
rect 916 -584 1052 -420
rect 1106 -586 1176 -420
rect 916 -1104 1052 -1030
rect 1106 -1104 1176 -1030
<< metal1 >>
rect 904 -264 1254 -194
rect 904 -408 1004 -264
rect 1046 -380 1112 -316
rect 904 -420 1052 -408
rect 904 -584 916 -420
rect 904 -598 1052 -584
rect 1106 -420 1184 -408
rect 1176 -586 1184 -420
rect 1106 -598 1184 -586
rect 1050 -784 1108 -634
rect 1030 -842 1040 -784
rect 1050 -990 1108 -842
rect 1136 -780 1184 -598
rect 1136 -786 1204 -780
rect 1136 -838 1146 -786
rect 1198 -838 1204 -786
rect 1136 -844 1204 -838
rect 1136 -1018 1184 -844
rect 904 -1030 1052 -1018
rect 904 -1104 916 -1030
rect 904 -1116 1052 -1104
rect 1106 -1030 1184 -1018
rect 1176 -1104 1184 -1030
rect 1106 -1116 1184 -1104
rect 904 -1252 1004 -1116
rect 1046 -1200 1112 -1144
rect 904 -1322 1254 -1252
<< via1 >>
rect 1040 -842 1108 -784
rect 1146 -838 1198 -786
<< metal2 >>
rect 1040 -784 1108 -774
rect 904 -842 1040 -784
rect 1136 -786 1290 -784
rect 1136 -838 1146 -786
rect 1198 -838 1290 -786
rect 1136 -842 1290 -838
rect 1040 -852 1108 -842
use sky130_fd_pr__nfet_01v8_4A3DHF  XM1
timestamp 1728411784
transform 1 0 1431 0 1 -1651
box -211 -255 211 255
use sky130_fd_pr__pfet_01v8_hvt_HVTLRR  XM2
timestamp 0
transform 1 0 1062 0 1 -1544
box -211 -309 211 309
<< labels >>
flabel metal2 1254 -842 1290 -784 0 FreeSans 256 0 0 0 Out
port 1 nsew
flabel metal2 904 -842 940 -784 0 FreeSans 256 0 0 0 In
port 2 nsew
flabel metal1 904 -264 1104 -194 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 904 -1322 1104 -1252 0 FreeSans 256 0 0 0 VSS
port 3 nsew
<< end >>
