* Extracted by KLayout with SKY130 LVS runset on : 05/11/2024 16:26

.SUBCKT RO_LVT_101St_x1 RON GND DUT_Gate RO DUT_Header OUT VDD DUT_Footer
+ Drain_Sense Drain\x20Force Out
M$1 VDD OUT \$241 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$5 VDD \$241 \$243 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$9 VDD \$243 \$245 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$13 VDD \$245 \$247 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$17 VDD \$247 \$249 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$21 VDD \$249 \$251 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$25 VDD \$251 \$253 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$29 VDD \$253 \$255 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$33 VDD \$255 \$257 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$37 VDD \$257 \$259 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$41 VDD \$259 \$261 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$45 VDD \$261 \$263 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$49 VDD \$263 \$265 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$53 VDD \$265 \$267 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$57 VDD \$267 \$269 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$61 VDD \$269 \$271 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$65 VDD \$271 \$273 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$69 VDD \$273 \$275 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$73 VDD \$275 \$277 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$77 VDD \$277 \$279 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$81 VDD \$279 \$281 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$85 VDD \$281 \$283 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$89 VDD \$283 \$285 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$93 VDD \$285 \$287 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$97 VDD \$287 \$289 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$101 VDD \$289 \$291 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$105 VDD \$291 \$293 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$109 VDD \$293 \$295 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$113 VDD \$295 \$297 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$117 VDD \$297 \$299 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$121 VDD \$299 \$301 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$125 VDD \$301 \$303 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$129 VDD \$303 \$305 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$133 VDD \$305 \$307 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$137 VDD \$307 \$309 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$141 VDD \$309 \$311 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$145 VDD \$311 \$313 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$149 VDD \$313 \$315 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$153 VDD \$315 \$317 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$157 VDD \$317 \$319 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$161 VDD \$319 \$321 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$165 VDD \$321 \$323 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$169 VDD \$323 \$325 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$173 VDD \$325 \$327 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$177 \$821 \$327 \$189 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$181 VDD RON \$821 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$221 \$822 \$189 \$194 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$225 VDD DUT_Footer \$822 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$265 \$194 RO Drain_Sense VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$269 \$194 RO Drain\x20Force VDD sky130_fd_pr__pfet_01v8_lvt L=350000
+ W=19000000 AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$273 \$823 \$194 \$195 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$277 VDD RON \$823 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=190000000
+ AS=2.92125e+13 AD=2.92125e+13 PS=207050000 PD=207050000
M$317 VDD \$1948 OUT VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$321 VDD \$1950 \$1948 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$325 VDD \$1952 \$1950 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$329 VDD \$1954 \$1952 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$333 VDD \$1956 \$1954 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$337 VDD \$1958 \$1956 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$341 VDD \$1960 \$1958 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$345 VDD \$1962 \$1960 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$349 VDD \$1964 \$1962 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$353 VDD \$1966 \$1964 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$357 VDD \$1968 \$1966 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$361 VDD \$1970 \$1968 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$365 VDD \$1972 \$1970 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$369 VDD \$1974 \$1972 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$373 VDD \$1976 \$1974 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$377 VDD \$1978 \$1976 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$381 VDD \$1980 \$1978 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$385 VDD \$1982 \$1980 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$389 VDD \$1984 \$1982 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$393 VDD \$1986 \$1984 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$397 VDD \$1988 \$1986 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$401 VDD \$1990 \$1988 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$405 VDD \$1992 \$1990 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$409 VDD \$1994 \$1992 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$413 VDD \$1996 \$1994 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$417 VDD \$1998 \$1996 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$421 VDD \$2000 \$1998 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$425 VDD \$2002 \$2000 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$429 VDD \$2004 \$2002 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$433 VDD \$2006 \$2004 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$437 VDD \$2008 \$2006 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$441 VDD \$2010 \$2008 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$445 VDD \$2012 \$2010 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$449 VDD \$2014 \$2012 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$453 VDD \$2016 \$2014 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$457 VDD \$2018 \$2016 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$461 VDD \$2020 \$2018 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$465 VDD \$2022 \$2020 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$469 VDD \$2024 \$2022 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$473 VDD \$2026 \$2024 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$477 VDD \$2028 \$2026 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$481 VDD \$2030 \$2028 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$485 VDD \$2032 \$2030 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$489 VDD \$1918 \$2032 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$493 \$1916 VDD \$1918 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$494 \$1917 VDD \$1918 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$495 VDD \$1921 \$1918 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$499 \$1919 VDD \$1921 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$500 \$1920 VDD \$1921 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$501 VDD \$1924 \$1921 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$505 \$1922 VDD \$1924 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$506 \$1923 VDD \$1924 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$507 VDD \$1927 \$1924 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$511 \$189 RO DUT_Gate VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$512 \$1925 VDD \$1927 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$513 \$189 RO \$193 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$514 \$1926 VDD \$1927 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$515 VDD \$1930 \$1927 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$519 \$1928 VDD \$1930 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$520 \$1929 VDD \$1930 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$521 VDD \$1933 \$1930 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$525 \$1931 VDD \$1933 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$526 \$1932 VDD \$1933 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$527 VDD \$1936 \$1933 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$531 \$1934 VDD \$1936 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$532 \$1935 VDD \$1936 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$533 VDD \$1939 \$1936 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$537 \$1937 VDD \$1939 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$538 \$1938 VDD \$1939 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$539 VDD \$1942 \$1939 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$543 \$1940 VDD \$1942 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$544 \$1941 VDD \$1942 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$545 VDD Out \$1942 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$549 \$1943 VDD Out VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$550 \$1944 VDD Out VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$551 VDD \$195 Out VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=19000000
+ AS=4.275e+12 AD=4.275e+12 PS=30300000 PD=30300000
M$555 \$195 VDD GND VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$556 \$195 VDD \$196 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$557 \$189 \$327 \$192 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$559 \$192 RO GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.26e+13 AD=1.26e+13 PS=96000000 PD=96000000
M$579 \$194 \$189 \$191 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$581 \$191 DUT_Header GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=42000000
+ AS=1.26e+13 AD=1.26e+13 PS=96000000 PD=96000000
M$601 \$194 RON Drain_Sense GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$603 \$194 RON Drain\x20Force GND sky130_fd_pr__nfet_01v8_lvt L=350000
+ W=4200000 AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$605 \$195 \$194 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$607 \$1916 GND \$1918 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$608 \$1917 GND \$1918 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$609 \$1918 \$1921 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$611 \$1919 GND \$1921 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$612 \$1920 GND \$1921 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$613 \$1921 \$1924 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$615 \$1922 GND \$1924 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$616 \$1923 GND \$1924 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$617 \$1924 \$1927 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$619 \$189 RON DUT_Gate GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$620 \$1925 GND \$1927 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$621 \$189 RON \$193 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$622 \$1926 GND \$1927 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$623 \$1927 \$1930 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$625 \$1928 GND \$1930 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$626 \$1929 GND \$1930 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$627 \$1930 \$1933 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$629 \$1931 GND \$1933 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$630 \$1932 GND \$1933 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$631 \$1933 \$1936 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$633 \$1934 GND \$1936 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$634 \$1935 GND \$1936 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$635 \$1936 \$1939 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$637 \$1937 GND \$1939 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$638 \$1938 GND \$1939 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$639 \$1939 \$1942 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$641 \$1940 GND \$1942 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$642 \$1941 GND \$1942 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$643 \$1942 Out GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$645 \$1943 GND Out GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$646 \$1944 GND Out GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$647 Out \$195 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$649 \$195 RON GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$650 \$195 RON \$196 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$651 \$241 OUT GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$653 OUT \$1948 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$655 \$243 \$241 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$657 \$1948 \$1950 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$659 \$245 \$243 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$661 \$1950 \$1952 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$663 \$247 \$245 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$665 \$1952 \$1954 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$667 \$249 \$247 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$669 \$1954 \$1956 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$671 \$251 \$249 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$673 \$1956 \$1958 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$675 \$253 \$251 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$677 \$1958 \$1960 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$679 \$255 \$253 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$681 \$1960 \$1962 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$683 \$257 \$255 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$685 \$1962 \$1964 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$687 \$259 \$257 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$689 \$1964 \$1966 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$691 \$261 \$259 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$693 \$1966 \$1968 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$695 \$263 \$261 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$697 \$1968 \$1970 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$699 \$265 \$263 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$701 \$1970 \$1972 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$703 \$267 \$265 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$705 \$1972 \$1974 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$707 \$269 \$267 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$709 \$1974 \$1976 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$711 \$271 \$269 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$713 \$1976 \$1978 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$715 \$273 \$271 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$717 \$1978 \$1980 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$719 \$275 \$273 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$721 \$1980 \$1982 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$723 \$277 \$275 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$725 \$1982 \$1984 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$727 \$279 \$277 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$729 \$1984 \$1986 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$731 \$281 \$279 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$733 \$1986 \$1988 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$735 \$283 \$281 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$737 \$1988 \$1990 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$739 \$285 \$283 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$741 \$1990 \$1992 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$743 \$287 \$285 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$745 \$1992 \$1994 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$747 \$289 \$287 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$749 \$1994 \$1996 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$751 \$291 \$289 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$753 \$1996 \$1998 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$755 \$293 \$291 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$757 \$1998 \$2000 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$759 \$295 \$293 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$761 \$2000 \$2002 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$763 \$297 \$295 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$765 \$2002 \$2004 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$767 \$299 \$297 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$769 \$2004 \$2006 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$771 \$301 \$299 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$773 \$2006 \$2008 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$775 \$303 \$301 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$777 \$2008 \$2010 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$779 \$305 \$303 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$781 \$2010 \$2012 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$783 \$307 \$305 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$785 \$2012 \$2014 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$787 \$309 \$307 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$789 \$2014 \$2016 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$791 \$311 \$309 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$793 \$2016 \$2018 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$795 \$313 \$311 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$797 \$2018 \$2020 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$799 \$315 \$313 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$801 \$2020 \$2022 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$803 \$317 \$315 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$805 \$2022 \$2024 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$807 \$319 \$317 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$809 \$2024 \$2026 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$811 \$321 \$319 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$813 \$2026 \$2028 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$815 \$323 \$321 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$817 \$2028 \$2030 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$819 \$325 \$323 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$821 \$2030 \$2032 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$823 \$327 \$325 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$825 \$2032 \$1918 GND GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=4200000
+ AS=1.26e+12 AD=1.26e+12 PS=9600000 PD=9600000
M$827 \$243 GND \$1012 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$828 \$243 GND \$1014 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$829 \$245 GND \$1016 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$830 \$245 GND \$1018 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$831 \$241 GND \$1008 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$832 \$241 GND \$1010 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$833 \$241 VDD \$1008 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$834 \$241 VDD \$1010 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$835 \$243 VDD \$1012 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$836 \$243 VDD \$1014 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$837 \$245 VDD \$1016 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$838 \$245 VDD \$1018 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$839 \$1950 VDD \$2952 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$840 \$1950 VDD \$2954 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$841 OUT VDD \$2944 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$842 OUT VDD \$2946 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$843 OUT GND \$2944 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$844 OUT GND \$2946 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$845 \$1950 GND \$2952 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$846 \$1950 GND \$2954 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$847 \$1948 GND \$2948 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$848 \$1948 GND \$2950 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$849 \$1948 VDD \$2948 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$850 \$1948 VDD \$2950 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$851 \$257 GND \$1040 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$852 \$257 GND \$1042 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$853 \$253 GND \$1032 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$854 \$253 GND \$1034 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$855 \$253 VDD \$1032 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$856 \$253 VDD \$1034 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$857 \$257 VDD \$1040 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$858 \$257 VDD \$1042 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$859 \$255 VDD \$1036 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$860 \$255 VDD \$1038 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$861 \$255 GND \$1036 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$862 \$255 GND \$1038 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$863 \$251 GND \$1028 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$864 \$251 GND \$1030 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$865 \$247 GND \$1020 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$866 \$247 GND \$1022 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$867 \$247 VDD \$1020 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$868 \$247 VDD \$1022 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$869 \$251 VDD \$1028 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$870 \$251 VDD \$1030 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$871 \$249 VDD \$1024 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$872 \$249 VDD \$1026 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$873 \$249 GND \$1024 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$874 \$249 GND \$1026 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$875 \$1956 VDD \$2964 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$876 \$1956 VDD \$2966 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$877 \$1954 VDD \$2960 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$878 \$1954 VDD \$2962 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$879 \$1952 GND \$2956 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$880 \$1952 GND \$2958 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$881 \$1954 GND \$2960 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$882 \$1954 GND \$2962 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$883 \$1956 GND \$2964 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$884 \$1956 GND \$2966 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$885 \$1962 VDD \$2976 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$886 \$1962 VDD \$2978 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$887 \$1960 VDD \$2972 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$888 \$1960 VDD \$2974 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$889 \$1960 GND \$2972 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$890 \$1960 GND \$2974 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$891 \$1962 GND \$2976 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$892 \$1962 GND \$2978 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$893 \$1958 GND \$2968 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$894 \$1958 GND \$2970 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$895 \$1958 VDD \$2968 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$896 \$1958 VDD \$2970 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$897 \$1952 VDD \$2956 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$898 \$1952 VDD \$2958 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$899 \$269 GND \$1064 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$900 \$269 GND \$1066 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$901 \$267 GND \$1060 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$902 \$267 GND \$1062 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$903 \$267 VDD \$1060 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$904 \$267 VDD \$1062 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$905 \$269 VDD \$1064 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$906 \$269 VDD \$1066 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$907 \$263 GND \$1052 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$908 \$263 GND \$1054 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$909 \$259 GND \$1044 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$910 \$259 GND \$1046 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$911 \$259 VDD \$1044 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$912 \$259 VDD \$1046 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$913 \$263 VDD \$1052 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$914 \$263 VDD \$1054 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$915 \$261 VDD \$1048 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$916 \$261 VDD \$1050 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$917 \$261 GND \$1048 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$918 \$261 GND \$1050 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$919 \$1968 VDD \$2988 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$920 \$1968 VDD \$2990 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$921 \$1966 VDD \$2984 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$922 \$1966 VDD \$2986 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$923 \$1966 GND \$2984 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$924 \$1966 GND \$2986 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$925 \$1970 GND \$2992 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$926 \$1970 GND \$2994 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$927 \$1968 GND \$2988 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$928 \$1968 GND \$2990 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$929 \$1976 VDD \$3004 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$930 \$1976 VDD \$3006 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$931 \$1972 VDD \$2996 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$932 \$1972 VDD \$2998 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$933 \$1972 GND \$2996 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$934 \$1972 GND \$2998 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$935 \$1976 GND \$3004 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$936 \$1976 GND \$3006 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$937 \$1974 GND \$3000 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$938 \$1974 GND \$3002 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$939 \$1974 VDD \$3000 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$940 \$1974 VDD \$3002 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$941 \$265 VDD \$1056 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$942 \$265 VDD \$1058 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$943 \$265 GND \$1056 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$944 \$265 GND \$1058 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$945 \$1970 VDD \$2992 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$946 \$1970 VDD \$2994 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$947 \$283 GND \$1092 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$948 \$283 GND \$1094 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$949 \$281 GND \$1088 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$950 \$281 GND \$1090 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$951 \$279 GND \$1084 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$952 \$279 GND \$1086 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$953 \$279 VDD \$1084 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$954 \$279 VDD \$1086 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$955 \$283 VDD \$1092 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$956 \$283 VDD \$1094 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$957 \$281 VDD \$1088 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$958 \$281 VDD \$1090 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$959 \$275 GND \$1076 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$960 \$275 GND \$1078 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$961 \$273 GND \$1072 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$962 \$273 GND \$1074 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$963 \$273 VDD \$1072 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$964 \$273 VDD \$1074 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$965 \$275 VDD \$1076 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$966 \$275 VDD \$1078 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$967 \$1982 VDD \$3016 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$968 \$1982 VDD \$3018 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$969 \$1978 VDD \$3008 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$970 \$1978 VDD \$3010 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$971 \$1978 GND \$3008 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$972 \$1978 GND \$3010 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$973 \$1982 GND \$3016 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$974 \$1982 GND \$3018 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$975 \$1980 GND \$3012 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$976 \$1980 GND \$3014 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$977 \$1980 VDD \$3012 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$978 \$1980 VDD \$3014 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$979 \$1988 VDD \$3028 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$980 \$1988 VDD \$3030 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$981 \$1984 VDD \$3020 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$982 \$1984 VDD \$3022 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$983 \$1984 GND \$3020 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$984 \$1984 GND \$3022 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$985 \$1988 GND \$3028 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$986 \$1988 GND \$3030 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$987 \$1986 GND \$3024 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$988 \$1986 GND \$3026 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$989 \$1986 VDD \$3024 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$990 \$1986 VDD \$3026 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$991 \$277 VDD \$1080 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$992 \$277 VDD \$1082 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$993 \$277 GND \$1080 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$994 \$277 GND \$1082 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$995 \$271 VDD \$1068 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$996 \$271 VDD \$1070 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$997 \$271 GND \$1068 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$998 \$271 GND \$1070 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$999 \$1964 GND \$2980 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1000 \$1964 GND \$2982 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1001 \$1964 VDD \$2980 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1002 \$1964 VDD \$2982 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1003 \$295 GND \$1116 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1004 \$295 GND \$1118 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1005 \$291 GND \$1108 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1006 \$291 GND \$1110 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1007 \$293 GND \$1112 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1008 \$293 GND \$1114 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1009 \$291 VDD \$1108 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1010 \$291 VDD \$1110 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1011 \$295 VDD \$1116 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1012 \$295 VDD \$1118 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1013 \$293 VDD \$1112 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1014 \$293 VDD \$1114 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1015 \$289 GND \$1104 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1016 \$289 GND \$1106 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1017 \$285 GND \$1096 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1018 \$285 GND \$1098 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1019 \$285 VDD \$1096 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1020 \$285 VDD \$1098 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1021 \$289 VDD \$1104 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1022 \$289 VDD \$1106 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1023 \$287 VDD \$1100 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1024 \$287 VDD \$1102 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1025 \$287 GND \$1100 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1026 \$287 GND \$1102 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1027 \$1994 VDD \$3040 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1028 \$1994 VDD \$3042 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1029 \$1992 VDD \$3036 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1030 \$1992 VDD \$3038 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1031 \$1990 VDD \$3032 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1032 \$1990 VDD \$3034 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1033 \$1990 GND \$3032 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1034 \$1990 GND \$3034 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1035 \$1992 GND \$3036 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1036 \$1992 GND \$3038 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1037 \$1994 GND \$3040 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1038 \$1994 GND \$3042 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1039 \$2000 VDD \$3052 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1040 \$2000 VDD \$3054 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1041 \$1998 VDD \$3048 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1042 \$1998 VDD \$3050 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1043 \$1998 GND \$3048 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1044 \$1998 GND \$3050 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1045 \$2000 GND \$3052 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1046 \$2000 GND \$3054 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1047 \$1996 GND \$3044 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1048 \$1996 GND \$3046 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1049 \$1996 VDD \$3044 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1050 \$1996 VDD \$3046 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1051 \$307 GND \$1140 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1052 \$307 GND \$1142 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1053 \$303 GND \$1132 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1054 \$303 GND \$1134 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1055 \$305 GND \$1136 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1056 \$305 GND \$1138 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1057 \$305 VDD \$1136 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1058 \$305 VDD \$1138 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1059 \$307 VDD \$1140 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1060 \$307 VDD \$1142 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1061 \$301 GND \$1128 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1062 \$301 GND \$1130 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1063 \$297 GND \$1120 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1064 \$297 GND \$1122 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1065 \$297 VDD \$1120 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1066 \$297 VDD \$1122 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1067 \$301 VDD \$1128 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1068 \$301 VDD \$1130 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1069 \$299 VDD \$1124 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1070 \$299 VDD \$1126 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1071 \$299 GND \$1124 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1072 \$299 GND \$1126 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1073 \$2006 VDD \$3064 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1074 \$2006 VDD \$3066 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1075 \$2004 VDD \$3060 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1076 \$2004 VDD \$3062 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1077 \$2004 GND \$3060 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1078 \$2004 GND \$3062 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1079 \$2006 GND \$3064 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1080 \$2006 GND \$3066 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1081 \$2014 VDD \$3080 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1082 \$2014 VDD \$3082 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1083 \$2010 VDD \$3072 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1084 \$2010 VDD \$3074 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1085 \$2010 GND \$3072 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1086 \$2010 GND \$3074 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1087 \$2014 GND \$3080 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1088 \$2014 GND \$3082 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1089 \$2012 GND \$3076 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1090 \$2012 GND \$3078 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1091 \$2012 VDD \$3076 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1092 \$2012 VDD \$3078 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1093 \$303 VDD \$1132 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1094 \$303 VDD \$1134 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1095 \$2008 GND \$3068 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1096 \$2008 GND \$3070 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1097 \$2008 VDD \$3068 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1098 \$2008 VDD \$3070 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1099 \$2002 GND \$3056 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1100 \$2002 GND \$3058 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1101 \$2002 VDD \$3056 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1102 \$2002 VDD \$3058 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1103 \$321 GND \$1168 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1104 \$321 GND \$1170 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1105 \$319 GND \$1164 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1106 \$319 GND \$1166 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1107 \$317 GND \$1160 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1108 \$317 GND \$1162 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1109 \$317 VDD \$1160 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1110 \$317 VDD \$1162 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1111 \$319 VDD \$1164 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1112 \$319 VDD \$1166 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1113 \$313 GND \$1152 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1114 \$313 GND \$1154 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1115 \$311 GND \$1148 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1116 \$311 GND \$1150 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1117 \$311 VDD \$1148 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1118 \$311 VDD \$1150 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1119 \$313 VDD \$1152 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1120 \$313 VDD \$1154 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1121 \$2020 VDD \$3092 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1122 \$2020 VDD \$3094 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1123 \$2016 VDD \$3084 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1124 \$2016 VDD \$3086 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1125 \$2016 GND \$3084 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1126 \$2016 GND \$3086 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1127 \$2020 GND \$3092 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1128 \$2020 GND \$3094 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1129 \$2018 GND \$3088 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1130 \$2018 GND \$3090 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1131 \$2018 VDD \$3088 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1132 \$2018 VDD \$3090 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1133 \$2026 VDD \$3104 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1134 \$2026 VDD \$3106 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1135 \$2022 VDD \$3096 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1136 \$2022 VDD \$3098 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1137 \$2022 GND \$3096 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1138 \$2022 GND \$3098 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1139 \$2026 GND \$3104 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1140 \$2026 GND \$3106 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1141 \$2024 GND \$3100 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1142 \$2024 GND \$3102 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1143 \$2024 VDD \$3100 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1144 \$2024 VDD \$3102 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1145 \$315 VDD \$1156 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1146 \$315 VDD \$1158 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1147 \$315 GND \$1156 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1148 \$315 GND \$1158 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1149 \$327 GND \$1180 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1150 \$327 GND \$1182 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1151 \$323 GND \$1172 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1152 \$323 GND \$1174 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1153 \$323 VDD \$1172 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1154 \$323 VDD \$1174 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1155 \$327 VDD \$1180 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1156 \$327 VDD \$1182 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1157 \$325 VDD \$1176 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1158 \$325 VDD \$1178 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1159 \$325 GND \$1176 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1160 \$325 GND \$1178 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1161 \$2032 VDD \$3116 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1162 \$2032 VDD \$3118 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1163 \$2030 VDD \$3112 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1164 \$2030 VDD \$3114 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1165 \$2028 VDD \$3108 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1166 \$2028 VDD \$3110 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1167 \$2028 GND \$3108 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1168 \$2028 GND \$3110 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1169 \$2030 GND \$3112 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1170 \$2030 GND \$3114 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1171 \$2032 GND \$3116 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1172 \$2032 GND \$3118 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1173 \$321 VDD \$1168 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1174 \$321 VDD \$1170 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1175 \$309 VDD \$1144 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1176 \$309 VDD \$1146 VDD sky130_fd_pr__pfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1177 \$309 GND \$1144 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
M$1178 \$309 GND \$1146 GND sky130_fd_pr__nfet_01v8_lvt L=350000 W=450000
+ AS=135000000000 AD=135000000000 PS=1500000 PD=1500000
.ENDS RO_LVT_101St_x1
