** sch_path: /foss/designs/RO_Aging_UNICASS/TB/13St_TB.sch
**.subckt 13St_TB
V1 VDD GND 1.8
V2 RO GND 1.8
V3 RON GND 0
V4 DUT_Header GND 1.8
V5 DUT_Footer GND 0
x2 VDD OUT OUT_B GND Buffer
x1 VDD GND DUT_Footer DUT_Header net1 net2 RO RON net3 OUT RO_LVT_13St_x1
x3 VDD OUT_Div OUT_B GND DIV
**** begin user architecture code

.tran 250n 1.1m
.ic V(OUT)=0.1
.save all

 .lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/Buffer/Buffer.sym # of pins=4
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/Buffer/Buffer.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/Buffer/Buffer.sch
.subckt Buffer VDD IN OUT GND
*.iopin VDD
*.iopin GND
*.iopin IN
*.iopin OUT
x1 VDD IN IN_NEG GND inv_LVT
x2 VDD IN_NEG OUT GND inv_LVT
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/RO_LVT_13St_x1/RO_LVT_13St_x1.sym # of pins=10
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/RO_LVT_13St_x1/RO_LVT_13St_x1.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/RO_LVT_13St_x1/RO_LVT_13St_x1.sch
.subckt RO_LVT_13St_x1 VDD GND DUT_Footer DUT_Header Drain_Sense Drain_Force RO RON DUT_Gate OUT
*.iopin DUT_Footer
*.iopin DUT_Header
*.iopin Drain_Sense
*.iopin Drain_Force
*.iopin RON
*.iopin RO
*.iopin DUT_Gate
*.iopin OUT
*.iopin GND
*.iopin VDD
x1[1] VDD GND A[7] A[8] rovcel2_LVT
x1[2] VDD GND A[6] A[7] rovcel2_LVT
x1[3] VDD GND A[5] A[6] rovcel2_LVT
x1[4] VDD GND A[4] A[5] rovcel2_LVT
x1[5] VDD GND A[3] A[4] rovcel2_LVT
x1[6] VDD GND A[2] A[3] rovcel2_LVT
x1[7] VDD GND A[1] A[2] rovcel2_LVT
x1[8] VDD GND OUT A[1] rovcel2_LVT
x2 VDD GND A[8] A[9] rovcel2_LVT
x6 VDD GND A[12] OUT rovcel2_LVT
x3 VDD GND RON A[9] A[10] RO DUT_Gate rovcel3_LVT
x4 VDD A[12] GND RON A[11] rovcel4_LVT
x1 VDD GND Drain_Sense DUT_Footer DUT_Header Drain_Force A[10] A[11] RON RO rovcel1_x1_LVT
.ends


* expanding   symbol:  DIV.sym # of pins=4
** sym_path: /foss/designs/RO_Aging_UNICASS/DIV/DIV.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/DIV.sch
.subckt DIV VDD OUT IN GND
*.iopin GND
*.iopin IN
*.iopin VDD
*.iopin OUT
x1 VDD A[0] A[0] net2 IN GND FF
* noconn #net2
x2 VDD A[1] A[1] net3 A[0] GND FF
* noconn #net3
x3[7] VDD OUT OUT net1 A[8] GND FF
x3[6] VDD A[8] A[8] net1 A[7] GND FF
x3[5] VDD A[7] A[7] net1 A[6] GND FF
x3[4] VDD A[6] A[6] net1 A[5] GND FF
x3[3] VDD A[5] A[5] net1 A[4] GND FF
x3[2] VDD A[4] A[4] net1 A[3] GND FF
x3[1] VDD A[3] A[3] net1 A[2] GND FF
x3[0] VDD A[2] A[2] net1 A[1] GND FF
* noconn #net1
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/inv_LVT/inv_LVT.sym # of pins=4
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/inv_LVT/inv_LVT.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/inv_LVT/inv_LVT.sch
.subckt inv_LVT VDD IN OUT GND
*.iopin VDD
*.iopin IN
*.iopin OUT
*.iopin GND
XM1 OUT IN GND GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/rovcel2_LVT/rovcel2_LVT.sym # of pins=4
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/rovcel2_LVT/rovcel2_LVT.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/rovcel2_LVT/rovcel2_LVT.sch
.subckt rovcel2_LVT VDD GND IN OUT
*.iopin OUT
*.iopin IN
*.iopin VDD
*.iopin GND
* noconn #net1
* noconn #net2
x1 VDD IN OUT GND inv_LVT
x2 VDD OUT net1 GND GND VDD passgate_LVT
x3 VDD OUT net2 GND GND VDD passgate_LVT
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/rovcel3_LVT/rovcel3_LVT.sym # of pins=7
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/rovcel3_LVT/rovcel3_LVT.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/rovcel3_LVT/rovcel3_LVT.sch
.subckt rovcel3_LVT VDD GND RON IN OUT RO DUT_Gate
*.iopin OUT
*.iopin DUT_Gate
*.iopin RON
*.iopin RO
*.iopin IN
*.iopin VDD
*.iopin GND
XM0 net2 RO GND GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20
XM1 OUT IN net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM2 OUT IN net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM3 net1 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=40 m=40
* noconn #net3
x2 RO OUT net3 RON GND VDD passgate_LVT
x3 RO OUT DUT_Gate RON GND VDD passgate_LVT
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/rovcel4_LVT/rovcel4_LVT.sym # of pins=5
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/rovcel4_LVT/rovcel4_LVT.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/rovcel4_LVT/rovcel4_LVT.sch
.subckt rovcel4_LVT VDD OUT GND RON IN
*.iopin OUT
*.iopin RON
*.iopin IN
*.iopin GND
*.iopin VDD
XM1 OUT IN GND GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM2 OUT IN net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM3 net1 RON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=40 m=40
* noconn #net2
x2 VDD OUT net2 RON GND VDD passgate_LVT
x3 VDD OUT GND RON GND VDD passgate_LVT
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/rovcel1_x1_LVT/rovcel1_x1_LVT.sym # of pins=10
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/rovcel1_x1_LVT/rovcel1_x1_LVT.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/rovcel1_x1_LVT/rovcel1_x1_LVT.sch
.subckt rovcel1_x1_LVT VDD GND Drain_Sense DUT_Footer DUT_Header Drain_Force IN OUT RON RO
*.iopin OUT
*.iopin Drain_Force
*.iopin DUT_Footer
*.iopin DUT_Header
*.iopin IN
*.iopin Drain_Sense
*.iopin VDD
*.iopin GND
*.iopin RO
*.iopin RON
XM0 net2 DUT_Header GND GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=20 m=20
XM1 OUT IN net2 GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=2.1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM2 OUT IN net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
XM3 net1 DUT_Footer VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=40 m=40
XM4 Drain_Force RON OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 Drain_Sense RON OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.42 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 Drain_Sense RO OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Drain_Force RO OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1.9 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/DIV/FF/FF.sym # of pins=6
** sym_path: /foss/designs/RO_Aging_UNICASS/DIV/FF/FF.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/FF/FF.sch
.subckt FF VDD D Q_N Q CLK GND
*.iopin GND
*.iopin CLK
*.iopin VDD
*.iopin Q
*.iopin Q_N
*.iopin D
x1 CLKN VDD net1 D GND CLK passgate_DIV
x2 VDD net2 net1 GND inv_DIV
x3 CLK VDD net1 net4 GND CLKN passgate_DIV
x4 VDD net4 net2 GND inv_DIV
x5 CLK VDD net3 net2 GND CLKN passgate_DIV
x6 VDD net5 net3 GND inv_DIV
x7 CLKN VDD net3 Q_N GND CLK passgate_DIV
x8 VDD Q Q_N GND inv_DIV
x10 VDD CLKN CLK GND inv_DIV
x9 VDD Q_N net5 GND inv_DIV
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/LVT/passgate_LVT/passgate_LVT.sym # of pins=6
** sym_path: /foss/designs/RO_Aging_UNICASS/LVT/passgate_LVT/passgate_LVT.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/LVT/passgate_LVT/passgate_LVT.sch
.subckt passgate_LVT CLKN IN OUT CLK GND VDD
*.iopin CLKN
*.iopin CLK
*.iopin IN
*.iopin OUT
*.iopin VDD
*.iopin GND
XM3 IN CLK OUT GND sky130_fd_pr__nfet_01v8_lvt L=0.35 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 IN CLKN OUT VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/DIV/passgate_DIV/passgate_DIV.sym # of pins=6
** sym_path: /foss/designs/RO_Aging_UNICASS/DIV/passgate_DIV/passgate_DIV.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/passgate_DIV/passgate_DIV.sch
.subckt passgate_DIV CLKN VDD OUT IN GND CLK
*.iopin VDD
*.iopin OUT
*.iopin GND
*.iopin IN
*.iopin CLKN
*.iopin CLK
XM3 IN CLK OUT GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 IN CLKN OUT VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/RO_Aging_UNICASS/DIV/inv_DIV/inv_DIV.sym # of pins=4
** sym_path: /foss/designs/RO_Aging_UNICASS/DIV/inv_DIV/inv_DIV.sym
** sch_path: /foss/designs/RO_Aging_UNICASS/DIV/inv_DIV/inv_DIV.sch
.subckt inv_DIV VDD OUT IN GND
*.iopin VDD
*.iopin OUT
*.iopin GND
*.iopin IN
XM3 OUT IN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
